# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

# High density, single height
SITE unithd
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.46 BY 2.72 ;
END unithd

# High density, double height
SITE unithddbl
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

LAYER nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END pwell

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.46 0.34 ;
  OFFSET 0.23 0.17 ;

  WIDTH 0.17 ;          # LI 1
  # SPACING  0.17 ;     # LI 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.17 ;
  AREA 0.0561 ;         # LI 6
  THICKNESS 0.1 ;
  EDGECAPACITANCE 40.697E-6 ;
  CAPACITANCE CPERSQDIST 36.9866E-6 ;
  RESISTANCE RPERSQ 12.2 ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 75 ) ( 0.0125 75 ) ( 0.0225 85.125 ) ( 22.5 10200 ) ) ;
END li1

LAYER mcon
  TYPE CUT ;

  WIDTH 0.17 ;                # Mcon 1
  SPACING 0.19 ;              # Mcon 2
  ENCLOSURE BELOW 0 0 ;       # Mcon 4
  ENCLOSURE ABOVE 0.03 0.06 ; # Met1 4 / Met1 5

  ANTENNADIFFAREARATIO PWL ( ( 0 3 ) ( 0.0125 3 ) ( 0.0225 3.405 ) ( 22.5 408 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.36 ; # mA per via Iavg_max at Tj = 90oC

END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 0.34 ;
  OFFSET 0.17 ;

  WIDTH 0.14 ;                     # Met1 1
  # SPACING 0.14 ;                 # Met1 2
  # SPACING 0.28 RANGE 3.001 100 ; # Met1 3b
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.14
     WIDTH 3 0.28 ;
  AREA 0.083 ;                     # Met1 6
  THICKNESS 0.35 ;
  MINENCLOSEDAREA 0.14 ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  EDGECAPACITANCE 40.567E-6 ;
  CAPACITANCE CPERSQDIST 25.7784E-6 ;
  DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;

  RESISTANCE RPERSQ 0.125 ;
END met1

LAYER via
  TYPE CUT ;
  WIDTH 0.15 ;                  # Via 1a
  SPACING 0.17 ;                # Via 2
  ENCLOSURE BELOW 0.055 0.085 ; # Via 4a / Via 5a
  ENCLOSURE ABOVE 0.055 0.085 ; # Met2 4 / Met2 5

  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.29 ; # mA per via Iavg_max at Tj = 90oC
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.46 ;
  OFFSET 0.23 ;

  WIDTH 0.14 ;                        # Met2 1
  # SPACING  0.14 ;                   # Met2 2
  # SPACING  0.28 RANGE 3.001 100 ;   # Met2 3b
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.14
     WIDTH 3 0.28 ;
  AREA 0.0676 ;                       # Met2 6
  THICKNESS 0.35 ;
  MINENCLOSEDAREA 0.14 ;

  EDGECAPACITANCE 37.759E-6 ;
  CAPACITANCE CPERSQDIST 16.9423E-6 ;
  RESISTANCE RPERSQ 0.125 ;
  DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;
END met2

# ******** Layer via2, type routing, number 44 **************
LAYER via2
  TYPE CUT ;
  WIDTH 0.2 ;                   # Via2 1
  SPACING 0.2 ;                 # Via2 2
  ENCLOSURE BELOW 0.04 0.085 ;  # Via2 4
  ENCLOSURE ABOVE 0.065 0.065 ; # Met3 4
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 0.68 ;
  OFFSET 0.34 ;

  WIDTH 0.3 ;              # Met3 1
  # SPACING 0.3 ;          # Met3 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.3
     WIDTH 3 0.4 ;
  AREA 0.24 ;              # Met3 6
  THICKNESS 0.8 ;

  EDGECAPACITANCE 40.989E-6 ;
  CAPACITANCE CPERSQDIST 12.3729E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;
END met3

LAYER via3
  TYPE CUT ;
  WIDTH 0.2 ;                   # Via3 1
  SPACING 0.2 ;                 # Via3 2
  ENCLOSURE BELOW 0.06 0.09 ;   # Via3 4 / Via3 5
  ENCLOSURE ABOVE 0.065 0.065 ; # Met4 3
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.92 ;
  OFFSET 0.46 ;

  WIDTH 0.3 ;             # Met4 1
  # SPACING  0.3 ;             # Met4 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.3
     WIDTH 3 0.4 ;
  AREA 0.24 ;            # Met4 4a

  THICKNESS 0.8 ;

  EDGECAPACITANCE 36.676E-6 ;
  CAPACITANCE CPERSQDIST 8.41537E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;
END met4

LAYER via4
  TYPE CUT ;

  WIDTH 0.8 ;                 # Via4 1
  SPACING 0.8 ;               # Via4 2
  ENCLOSURE BELOW 0.19 0.19 ; # Via4 4
  ENCLOSURE ABOVE 0.31 0.31 ; # Met5 3
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 2.49 ; # mA per via Iavg_max at Tj = 90oC
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 3.4 ;
  OFFSET 1.7 ;

  WIDTH 1.6 ;            # Met5 1
  #SPACING  1.6 ;        # Met5 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 1.6 ;
  AREA 4 ;               # Met5 4

  THICKNESS 1.2 ;

  EDGECAPACITANCE 38.851E-6 ;
  CAPACITANCE CPERSQDIST 6.32063E-6 ;
  RESISTANCE RPERSQ 0.0285 ;
  DCCURRENTDENSITY AVERAGE 10.17 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 22.34 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met5


### Routing via cells section   ###
# Plus via rule, metals are along the prefered direction
VIA L1M1_PR DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIARULE L1M1_PR GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.03 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR

# Plus via rule, metals are along the non prefered direction
VIA L1M1_PR_R DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIARULE L1M1_PR_R GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.03 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA L1M1_PR_M DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIARULE L1M1_PR_M GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.03 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA L1M1_PR_MR DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIARULE L1M1_PR_MR GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.03 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_MR

# Centered via rule, we really do not want to use it
VIA L1M1_PR_C DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIARULE L1M1_PR_C GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_C

# Plus via rule, metals are along the prefered direction
VIA M1M2_PR DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.13 0.16 0.13 ;
  LAYER met2 ;
  RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIARULE M1M2_PR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER met2 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR

# Plus via rule, metals are along the non prefered direction
VIA M1M2_PR_R DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.13 -0.16 0.13 0.16 ;
  LAYER met2 ;
  RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIARULE M1M2_PR_R GENERATE
  LAYER met1 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M1M2_PR_M DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.13 0.16 0.13 ;
  LAYER met2 ;
  RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIARULE M1M2_PR_M GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M1M2_PR_MR DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.13 -0.16 0.13 0.16 ;
  LAYER met2 ;
  RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIARULE M1M2_PR_MR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_MR

# Centered via rule, we really do not want to use it
VIA M1M2_PR_C DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.16 0.16 0.16 ;
  LAYER met2 ;
  RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIARULE M1M2_PR_C GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_C

# Plus via rule, metals are along the prefered direction
VIA M2M3_PR DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.14 -0.185 0.14 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIARULE M2M3_PR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.04 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR

# Plus via rule, metals are along the non prefered direction
VIA M2M3_PR_R DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.14 0.185 0.14 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIARULE M2M3_PR_R GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.04 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M2M3_PR_M DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.14 -0.185 0.14 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIARULE M2M3_PR_M GENERATE
  LAYER met2 ;
  ENCLOSURE 0.04 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M2M3_PR_MR DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.14 0.185 0.14 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIARULE M2M3_PR_MR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.04 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_MR

# Centered via rule, we really do not want to use it
VIA M2M3_PR_C DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.185 0.185 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIARULE M2M3_PR_C GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_C

# Plus via rule, metals are along the prefered direction
VIA M3M4_PR DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.16 0.19 0.16 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIARULE M3M4_PR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.06 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR

# Plus via rule, metals are along the non prefered direction
VIA M3M4_PR_R DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.16 -0.19 0.16 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIARULE M3M4_PR_R GENERATE
  LAYER met3 ;
  ENCLOSURE 0.06 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M3M4_PR_M DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.16 0.19 0.16 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIARULE M3M4_PR_M GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.06 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M3M4_PR_MR DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.16 -0.19 0.16 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIARULE M3M4_PR_MR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.06 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_MR

# Centered via rule, we really do not want to use it
VIA M3M4_PR_C DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.19 0.19 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIARULE M3M4_PR_C GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_C

# Plus via rule, metals are along the prefered direction
VIA M4M5_PR DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIARULE M4M5_PR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR

# Plus via rule, metals are along the non prefered direction
VIA M4M5_PR_R DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIARULE M4M5_PR_R GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M4M5_PR_M DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIARULE M4M5_PR_M GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M4M5_PR_MR DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIARULE M4M5_PR_MR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_MR

# Centered via rule, we really do not want to use it
VIA M4M5_PR_C DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

VIARULE M4M5_PR_C GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_C
###  end of single via cells   ###


MACRO sky130_ef_sc_hd__fakediode_2
  CLASS CORE SPACER ;
  FOREIGN sky130_ef_sc_hd__fakediode_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.920000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DIODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.835000 2.465000 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.920000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.110000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.920000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.920000 0.085000 ;
      RECT 0.000000  2.635000 0.920000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
  END
END sky130_ef_sc_hd__fakediode_2
MACRO sky130_ef_sc_hd__fill_8
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.680000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.680000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
  END
END sky130_ef_sc_hd__fill_8
MACRO sky130_ef_sc_hd__decap_12
  CLASS BLOCK ;
  FOREIGN sky130_ef_sc_hd__decap_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 1.670 0.630 2.010 1.460 ;
        RECT 0.085 0.085 5.430 0.630 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INPUT ;
    PORT
      LAYER pwell ;
        RECT 0.080 -0.130 0.360 0.150 ;
    END
  END VNB
  PIN VPB
    DIRECTION INPUT ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.085 2.200 5.430 2.635 ;
        RECT 3.490 0.950 3.840 2.200 ;
      LAYER mcon ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
END sky130_ef_sc_hd__decap_12
MACRO sky130_ef_sc_hd__fill_12
  CLASS CORE ;
  FOREIGN sky130_ef_sc_hd__fill_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 2.935 -0.060 3.045 0.060 ;
        RECT 4.755 -0.050 4.915 0.060 ;
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.085 1.545 2.675 2.635 ;
        RECT 0.085 0.855 1.295 1.375 ;
        RECT 1.465 1.025 2.675 1.545 ;
        RECT 0.085 0.085 2.675 0.855 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
        RECT 0.000 -0.240 5.520 0.240 ;
  END
END sky130_ef_sc_hd__fill_12
MACRO sky130_fd_sc_hd__a2bb2o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.910000 0.995000 1.240000 1.615000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.410000 0.995000 1.700000 1.375000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.280000 0.765000 3.540000 1.655000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.600000 1.355000 3.080000 1.655000 ;
        RECT 2.820000 0.765000 3.080000 1.355000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.345000 0.810000 ;
        RECT 0.085000 0.810000 0.260000 1.525000 ;
        RECT 0.085000 1.525000 0.345000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.430000  0.995000 0.685000 1.325000 ;
      RECT 0.515000  0.085000 0.945000 0.530000 ;
      RECT 0.515000  1.325000 0.685000 1.805000 ;
      RECT 0.515000  1.805000 1.275000 1.975000 ;
      RECT 0.515000  2.235000 0.845000 2.635000 ;
      RECT 1.105000  1.975000 1.275000 2.200000 ;
      RECT 1.105000  2.200000 2.245000 2.370000 ;
      RECT 1.180000  0.255000 1.350000 0.655000 ;
      RECT 1.180000  0.655000 2.060000 0.825000 ;
      RECT 1.520000  0.085000 2.240000 0.485000 ;
      RECT 1.540000  1.545000 2.060000 1.715000 ;
      RECT 1.540000  1.715000 1.710000 1.905000 ;
      RECT 1.890000  0.825000 2.060000 1.545000 ;
      RECT 1.990000  1.895000 2.400000 2.065000 ;
      RECT 1.990000  2.065000 2.245000 2.200000 ;
      RECT 1.990000  2.370000 2.245000 2.465000 ;
      RECT 2.230000  0.700000 2.580000 0.870000 ;
      RECT 2.230000  0.870000 2.400000 1.895000 ;
      RECT 2.410000  0.255000 2.580000 0.700000 ;
      RECT 2.415000  2.255000 2.745000 2.425000 ;
      RECT 2.575000  1.835000 3.515000 2.005000 ;
      RECT 2.575000  2.005000 2.745000 2.255000 ;
      RECT 2.915000  2.175000 3.165000 2.635000 ;
      RECT 3.155000  0.085000 3.555000 0.595000 ;
      RECT 3.335000  2.005000 3.515000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a2bb2o_1
MACRO sky130_fd_sc_hd__a2bb2o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.345000 0.995000 1.675000 1.615000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.845000 0.995000 2.135000 1.375000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.730000 0.765000 3.990000 1.655000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.050000 1.355000 3.530000 1.655000 ;
        RECT 3.270000 0.765000 3.530000 1.355000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 0.255000 0.780000 0.810000 ;
        RECT 0.525000 0.810000 0.695000 1.525000 ;
        RECT 0.525000 1.525000 0.780000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.125000 -0.085000 0.295000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.185000  0.085000 0.355000 0.930000 ;
      RECT 0.185000  1.445000 0.355000 2.635000 ;
      RECT 0.865000  0.995000 1.120000 1.325000 ;
      RECT 0.950000  0.085000 1.380000 0.530000 ;
      RECT 0.950000  1.325000 1.120000 1.805000 ;
      RECT 0.950000  1.805000 1.710000 1.975000 ;
      RECT 0.950000  2.235000 1.280000 2.635000 ;
      RECT 1.540000  1.975000 1.710000 2.200000 ;
      RECT 1.540000  2.200000 2.670000 2.370000 ;
      RECT 1.615000  0.255000 1.785000 0.655000 ;
      RECT 1.615000  0.655000 2.510000 0.825000 ;
      RECT 1.955000  0.085000 2.690000 0.485000 ;
      RECT 1.975000  1.545000 2.510000 1.715000 ;
      RECT 1.975000  1.715000 2.145000 1.905000 ;
      RECT 2.340000  0.825000 2.510000 1.545000 ;
      RECT 2.440000  1.895000 2.850000 2.065000 ;
      RECT 2.440000  2.065000 2.670000 2.200000 ;
      RECT 2.500000  2.370000 2.670000 2.465000 ;
      RECT 2.680000  0.700000 3.030000 0.870000 ;
      RECT 2.680000  0.870000 2.850000 1.895000 ;
      RECT 2.860000  0.255000 3.030000 0.700000 ;
      RECT 2.875000  2.255000 3.205000 2.425000 ;
      RECT 3.035000  1.835000 3.965000 2.005000 ;
      RECT 3.035000  2.005000 3.205000 2.255000 ;
      RECT 3.375000  2.175000 3.625000 2.635000 ;
      RECT 3.605000  0.085000 4.005000 0.595000 ;
      RECT 3.795000  2.005000 3.965000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__a2bb2o_2
MACRO sky130_fd_sc_hd__a2bb2o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 1.075000 3.645000 1.325000 ;
        RECT 3.475000 1.325000 3.645000 1.445000 ;
        RECT 3.475000 1.445000 4.965000 1.615000 ;
        RECT 4.605000 1.075000 4.965000 1.445000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 1.075000 4.435000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.575000 1.445000 ;
        RECT 0.085000 1.445000 1.685000 1.615000 ;
        RECT 1.515000 1.075000 1.895000 1.245000 ;
        RECT 1.515000 1.245000 1.685000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 1.075000 1.345000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235000 0.275000 5.565000 0.725000 ;
        RECT 5.235000 0.725000 6.920000 0.905000 ;
        RECT 5.275000 1.785000 6.365000 1.955000 ;
        RECT 5.275000 1.955000 5.525000 2.465000 ;
        RECT 6.075000 0.275000 6.405000 0.725000 ;
        RECT 6.115000 1.415000 6.920000 1.655000 ;
        RECT 6.115000 1.655000 6.365000 1.785000 ;
        RECT 6.115000 1.955000 6.365000 2.465000 ;
        RECT 6.610000 0.905000 6.920000 1.415000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.135000  1.785000 2.065000 1.955000 ;
      RECT 0.135000  1.955000 0.385000 2.465000 ;
      RECT 0.175000  0.085000 0.345000 0.895000 ;
      RECT 0.515000  0.255000 1.685000 0.475000 ;
      RECT 0.515000  0.475000 0.765000 0.905000 ;
      RECT 0.555000  2.125000 0.805000 2.635000 ;
      RECT 0.935000  0.645000 1.270000 0.735000 ;
      RECT 0.935000  0.735000 2.525000 0.905000 ;
      RECT 0.975000  1.955000 1.225000 2.465000 ;
      RECT 1.395000  2.125000 1.645000 2.635000 ;
      RECT 1.815000  1.955000 2.065000 2.295000 ;
      RECT 1.815000  2.295000 2.905000 2.465000 ;
      RECT 1.855000  0.085000 2.025000 0.555000 ;
      RECT 1.855000  1.455000 2.065000 1.785000 ;
      RECT 2.195000  0.255000 2.525000 0.735000 ;
      RECT 2.235000  0.905000 2.445000 1.415000 ;
      RECT 2.235000  1.415000 2.620000 1.965000 ;
      RECT 2.235000  1.965000 2.485000 2.125000 ;
      RECT 2.615000  1.075000 3.145000 1.245000 ;
      RECT 2.655000  2.135000 2.905000 2.295000 ;
      RECT 2.695000  0.085000 3.385000 0.555000 ;
      RECT 2.955000  0.725000 4.725000 0.905000 ;
      RECT 2.955000  0.905000 3.145000 1.075000 ;
      RECT 2.955000  1.245000 3.145000 1.495000 ;
      RECT 2.955000  1.495000 3.305000 1.665000 ;
      RECT 3.135000  1.665000 3.305000 1.785000 ;
      RECT 3.135000  1.785000 4.265000 1.965000 ;
      RECT 3.175000  2.135000 3.425000 2.635000 ;
      RECT 3.555000  0.255000 3.885000 0.725000 ;
      RECT 3.595000  2.135000 3.845000 2.295000 ;
      RECT 3.595000  2.295000 4.685000 2.465000 ;
      RECT 4.015000  1.965000 4.265000 2.125000 ;
      RECT 4.055000  0.085000 4.225000 0.555000 ;
      RECT 4.395000  0.255000 4.725000 0.725000 ;
      RECT 4.435000  1.785000 4.685000 2.295000 ;
      RECT 4.855000  1.795000 5.105000 2.635000 ;
      RECT 4.895000  0.085000 5.065000 0.895000 ;
      RECT 5.135000  1.075000 6.440000 1.245000 ;
      RECT 5.135000  1.245000 5.460000 1.615000 ;
      RECT 5.695000  2.165000 5.945000 2.635000 ;
      RECT 5.735000  0.085000 5.905000 0.555000 ;
      RECT 6.535000  1.825000 6.785000 2.635000 ;
      RECT 6.575000  0.085000 6.745000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.450000  1.445000 2.620000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.230000  1.445000 5.400000 1.615000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
    LAYER met1 ;
      RECT 2.390000 1.415000 2.680000 1.460000 ;
      RECT 2.390000 1.460000 5.460000 1.600000 ;
      RECT 2.390000 1.600000 2.680000 1.645000 ;
      RECT 5.170000 1.415000 5.460000 1.460000 ;
      RECT 5.170000 1.600000 5.460000 1.645000 ;
  END
END sky130_fd_sc_hd__a2bb2o_4
MACRO sky130_fd_sc_hd__a2bb2oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.995000 0.520000 1.615000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.725000 1.010000 1.240000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.780000 0.995000 3.070000 1.615000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.245000 0.995000 2.610000 1.615000 ;
        RECT 2.440000 0.425000 2.610000 0.995000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.515500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.420000 1.785000 1.945000 1.955000 ;
        RECT 1.420000 1.955000 1.785000 2.465000 ;
        RECT 1.775000 0.255000 2.205000 0.825000 ;
        RECT 1.775000 0.825000 1.945000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.825000 ;
      RECT 0.095000  1.805000 0.425000 2.635000 ;
      RECT 0.595000  0.255000 0.765000 0.660000 ;
      RECT 0.595000  0.660000 1.580000 0.830000 ;
      RECT 0.875000  1.445000 1.580000 1.615000 ;
      RECT 0.875000  1.615000 1.205000 2.465000 ;
      RECT 0.935000  0.085000 1.605000 0.490000 ;
      RECT 1.410000  0.830000 1.580000 1.445000 ;
      RECT 1.955000  2.235000 2.285000 2.465000 ;
      RECT 2.115000  1.785000 3.130000 1.955000 ;
      RECT 2.115000  1.955000 2.285000 2.235000 ;
      RECT 2.455000  2.135000 2.705000 2.635000 ;
      RECT 2.795000  0.085000 3.125000 0.825000 ;
      RECT 2.875000  1.955000 3.130000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a2bb2oi_1
MACRO sky130_fd_sc_hd__a2bb2oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.310000 1.075000 4.205000 1.275000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.455000 1.075000 5.435000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.710000 1.445000 ;
        RECT 0.085000 1.445000 2.030000 1.615000 ;
        RECT 1.700000 1.075000 2.030000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.940000 1.075000 1.480000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 0.645000 1.400000 0.725000 ;
        RECT 1.070000 0.725000 2.660000 0.905000 ;
        RECT 2.330000 0.255000 2.660000 0.725000 ;
        RECT 2.370000 0.905000 2.660000 1.660000 ;
        RECT 2.370000 1.660000 2.620000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.270000  1.785000 2.200000 1.955000 ;
      RECT 0.270000  1.955000 0.520000 2.465000 ;
      RECT 0.310000  0.085000 0.480000 0.895000 ;
      RECT 0.650000  0.255000 1.820000 0.475000 ;
      RECT 0.650000  0.475000 0.900000 0.895000 ;
      RECT 0.690000  2.135000 0.940000 2.635000 ;
      RECT 1.110000  1.955000 1.360000 2.465000 ;
      RECT 1.530000  2.135000 1.780000 2.635000 ;
      RECT 1.950000  1.955000 2.200000 2.295000 ;
      RECT 1.950000  2.295000 3.040000 2.465000 ;
      RECT 1.990000  0.085000 2.160000 0.555000 ;
      RECT 2.790000  1.795000 3.040000 2.295000 ;
      RECT 2.830000  0.085000 3.520000 0.555000 ;
      RECT 2.830000  0.995000 3.120000 1.325000 ;
      RECT 2.950000  0.725000 4.860000 0.905000 ;
      RECT 2.950000  0.905000 3.120000 0.995000 ;
      RECT 2.950000  1.325000 3.120000 1.445000 ;
      RECT 2.950000  1.445000 4.820000 1.615000 ;
      RECT 3.310000  1.785000 4.400000 1.965000 ;
      RECT 3.310000  1.965000 3.560000 2.465000 ;
      RECT 3.690000  0.255000 4.020000 0.725000 ;
      RECT 3.730000  2.135000 3.980000 2.635000 ;
      RECT 4.150000  1.965000 4.400000 2.295000 ;
      RECT 4.150000  2.295000 5.240000 2.465000 ;
      RECT 4.190000  0.085000 4.360000 0.555000 ;
      RECT 4.530000  0.255000 4.860000 0.725000 ;
      RECT 4.570000  1.615000 4.820000 2.125000 ;
      RECT 4.990000  1.455000 5.240000 2.295000 ;
      RECT 5.030000  0.085000 5.200000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__a2bb2oi_2
MACRO sky130_fd_sc_hd__a2bb2oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.945000 1.075000 7.320000 1.275000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.595000 1.075000 9.045000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.075000 1.555000 1.285000 ;
        RECT 1.385000 1.285000 1.555000 1.445000 ;
        RECT 1.385000 1.445000 3.575000 1.615000 ;
        RECT 3.245000 1.075000 3.575000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.725000 1.075000 3.075000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775000 0.645000 2.995000 0.725000 ;
        RECT 1.775000 0.725000 5.045000 0.905000 ;
        RECT 3.745000 0.905000 3.915000 1.415000 ;
        RECT 3.745000 1.415000 4.965000 1.615000 ;
        RECT 3.875000 0.275000 4.205000 0.725000 ;
        RECT 3.915000 1.615000 4.165000 2.125000 ;
        RECT 4.715000 0.275000 5.045000 0.725000 ;
        RECT 4.745000 1.615000 4.965000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.085000  1.455000 1.215000 1.625000 ;
      RECT 0.085000  1.625000 0.425000 2.465000 ;
      RECT 0.175000  0.085000 0.345000 0.895000 ;
      RECT 0.515000  0.255000 0.845000 0.725000 ;
      RECT 0.515000  0.725000 1.605000 0.905000 ;
      RECT 0.595000  1.795000 0.805000 2.635000 ;
      RECT 0.975000  1.625000 1.215000 1.795000 ;
      RECT 0.975000  1.795000 3.745000 1.965000 ;
      RECT 0.975000  1.965000 1.215000 2.465000 ;
      RECT 1.015000  0.085000 1.185000 0.555000 ;
      RECT 1.355000  0.255000 3.365000 0.475000 ;
      RECT 1.355000  0.475000 1.605000 0.725000 ;
      RECT 1.395000  2.135000 1.645000 2.635000 ;
      RECT 1.815000  1.965000 2.065000 2.465000 ;
      RECT 2.235000  2.135000 2.485000 2.635000 ;
      RECT 2.655000  1.965000 2.905000 2.465000 ;
      RECT 3.075000  2.135000 3.325000 2.635000 ;
      RECT 3.495000  1.965000 3.745000 2.295000 ;
      RECT 3.495000  2.295000 5.465000 2.465000 ;
      RECT 3.535000  0.085000 3.705000 0.555000 ;
      RECT 4.085000  1.075000 5.725000 1.245000 ;
      RECT 4.335000  1.795000 4.575000 2.295000 ;
      RECT 4.375000  0.085000 4.545000 0.555000 ;
      RECT 5.135000  1.455000 5.465000 2.295000 ;
      RECT 5.215000  0.085000 5.905000 0.555000 ;
      RECT 5.555000  0.735000 9.575000 0.905000 ;
      RECT 5.555000  0.905000 5.725000 1.075000 ;
      RECT 5.655000  1.455000 7.625000 1.625000 ;
      RECT 5.655000  1.625000 5.985000 2.465000 ;
      RECT 6.075000  0.255000 6.405000 0.725000 ;
      RECT 6.075000  0.725000 8.925000 0.735000 ;
      RECT 6.155000  1.795000 6.365000 2.635000 ;
      RECT 6.540000  1.625000 6.780000 2.465000 ;
      RECT 6.575000  0.085000 6.745000 0.555000 ;
      RECT 6.915000  0.255000 7.245000 0.725000 ;
      RECT 6.955000  1.795000 7.205000 2.635000 ;
      RECT 7.375000  1.625000 7.625000 2.295000 ;
      RECT 7.375000  2.295000 9.310000 2.465000 ;
      RECT 7.415000  0.085000 7.585000 0.555000 ;
      RECT 7.755000  0.255000 8.085000 0.725000 ;
      RECT 7.795000  1.455000 9.575000 1.625000 ;
      RECT 7.795000  1.625000 8.045000 2.125000 ;
      RECT 8.215000  1.795000 8.465000 2.295000 ;
      RECT 8.255000  0.085000 8.425000 0.555000 ;
      RECT 8.595000  0.255000 8.925000 0.725000 ;
      RECT 8.635000  1.625000 8.885000 2.125000 ;
      RECT 9.060000  1.795000 9.310000 2.295000 ;
      RECT 9.095000  0.085000 9.265000 0.555000 ;
      RECT 9.215000  0.905000 9.575000 1.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
END sky130_fd_sc_hd__a2bb2oi_4
MACRO sky130_fd_sc_hd__a21bo_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21bo_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.750000 0.995000 2.175000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.370000 0.995000 2.630000 1.615000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.325000 0.335000 1.665000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.300000 0.265000 3.580000 2.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.105000  1.845000 0.855000 2.045000 ;
      RECT 0.105000  2.045000 0.345000 2.435000 ;
      RECT 0.515000  0.265000 0.745000 1.165000 ;
      RECT 0.515000  1.165000 0.855000 1.845000 ;
      RECT 0.515000  2.225000 0.865000 2.635000 ;
      RECT 0.945000  0.085000 1.190000 0.865000 ;
      RECT 1.035000  1.045000 1.580000 1.345000 ;
      RECT 1.035000  1.345000 1.365000 2.455000 ;
      RECT 1.360000  0.265000 1.790000 0.625000 ;
      RECT 1.360000  0.625000 3.100000 0.815000 ;
      RECT 1.360000  0.815000 1.580000 1.045000 ;
      RECT 1.535000  1.785000 2.560000 1.985000 ;
      RECT 1.535000  1.985000 1.715000 2.455000 ;
      RECT 1.885000  2.155000 2.215000 2.635000 ;
      RECT 2.370000  0.085000 3.100000 0.455000 ;
      RECT 2.390000  1.985000 2.560000 2.455000 ;
      RECT 2.825000  1.495000 3.110000 2.635000 ;
      RECT 2.840000  0.815000 3.100000 1.325000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a21bo_1
MACRO sky130_fd_sc_hd__a21bo_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21bo_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.685000 0.995000 3.100000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.270000 0.995000 3.560000 1.615000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 1.035000 1.525000 1.325000 ;
        RECT 1.330000 0.995000 1.525000 1.035000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.715000 0.850000 0.885000 ;
        RECT 0.150000 0.885000 0.380000 1.835000 ;
        RECT 0.150000 1.835000 0.850000 2.005000 ;
        RECT 0.520000 0.315000 0.850000 0.715000 ;
        RECT 0.595000 2.005000 0.850000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.090000  0.085000 0.345000 0.545000 ;
      RECT 0.090000  2.255000 0.425000 2.635000 ;
      RECT 0.570000  1.075000 0.900000 1.495000 ;
      RECT 0.570000  1.495000 1.285000 1.665000 ;
      RECT 1.020000  0.085000 1.220000 0.865000 ;
      RECT 1.040000  2.275000 1.370000 2.635000 ;
      RECT 1.115000  1.665000 1.285000 1.895000 ;
      RECT 1.115000  1.895000 2.225000 2.105000 ;
      RECT 1.455000  0.655000 1.865000 0.825000 ;
      RECT 1.455000  1.555000 1.865000 1.725000 ;
      RECT 1.695000  0.825000 1.865000 0.995000 ;
      RECT 1.695000  0.995000 2.175000 1.325000 ;
      RECT 1.695000  1.325000 1.865000 1.555000 ;
      RECT 1.975000  0.085000 2.305000 0.465000 ;
      RECT 1.975000  2.105000 2.225000 2.465000 ;
      RECT 2.055000  1.505000 2.515000 1.675000 ;
      RECT 2.055000  1.675000 2.225000 1.895000 ;
      RECT 2.345000  0.635000 2.740000 0.825000 ;
      RECT 2.345000  0.825000 2.515000 1.505000 ;
      RECT 2.395000  1.845000 3.565000 2.015000 ;
      RECT 2.395000  2.015000 2.725000 2.465000 ;
      RECT 2.895000  2.185000 3.065000 2.635000 ;
      RECT 3.235000  0.085000 3.565000 0.825000 ;
      RECT 3.235000  2.015000 3.565000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a21bo_2
MACRO sky130_fd_sc_hd__a21bo_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21bo_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.590000 1.010000 4.955000 1.360000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.025000 1.010000 4.420000 1.275000 ;
        RECT 4.245000 1.275000 4.420000 1.595000 ;
        RECT 4.245000 1.595000 5.390000 1.765000 ;
        RECT 5.220000 1.055000 5.700000 1.290000 ;
        RECT 5.220000 1.290000 5.390000 1.595000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.500000 1.010000 0.830000 1.625000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 0.615000 2.340000 0.785000 ;
        RECT 1.000000 0.785000 1.235000 1.595000 ;
        RECT 1.000000 1.595000 2.410000 1.765000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.105000  0.255000 0.540000 0.840000 ;
      RECT 0.105000  0.840000 0.330000 1.795000 ;
      RECT 0.105000  1.795000 0.565000 1.935000 ;
      RECT 0.105000  1.935000 2.870000 2.105000 ;
      RECT 0.105000  2.105000 0.550000 2.465000 ;
      RECT 0.710000  0.085000 1.050000 0.445000 ;
      RECT 0.720000  2.275000 1.050000 2.635000 ;
      RECT 1.405000  0.995000 2.810000 1.185000 ;
      RECT 1.405000  1.185000 2.530000 1.325000 ;
      RECT 1.580000  0.085000 1.910000 0.445000 ;
      RECT 1.580000  2.275000 1.910000 2.635000 ;
      RECT 2.435000  2.275000 2.770000 2.635000 ;
      RECT 2.515000  0.085000 3.285000 0.445000 ;
      RECT 2.640000  0.615000 3.645000 0.670000 ;
      RECT 2.640000  0.670000 4.965000 0.785000 ;
      RECT 2.640000  0.785000 3.010000 0.800000 ;
      RECT 2.640000  0.800000 2.810000 0.995000 ;
      RECT 2.700000  1.355000 3.305000 1.525000 ;
      RECT 2.700000  1.525000 2.870000 1.935000 ;
      RECT 2.995000  0.995000 3.305000 1.355000 ;
      RECT 3.055000  1.695000 3.225000 2.210000 ;
      RECT 3.055000  2.210000 4.065000 2.380000 ;
      RECT 3.475000  0.255000 3.645000 0.615000 ;
      RECT 3.475000  0.785000 4.965000 0.840000 ;
      RECT 3.475000  0.840000 3.645000 1.805000 ;
      RECT 3.855000  0.085000 4.185000 0.445000 ;
      RECT 3.885000  1.445000 4.065000 1.935000 ;
      RECT 3.885000  1.935000 5.825000 2.105000 ;
      RECT 3.885000  2.105000 4.065000 2.210000 ;
      RECT 4.235000  2.275000 4.565000 2.635000 ;
      RECT 4.685000  0.405000 4.965000 0.670000 ;
      RECT 5.075000  2.275000 5.405000 2.635000 ;
      RECT 5.545000  0.085000 5.825000 0.885000 ;
      RECT 5.570000  1.460000 5.825000 1.935000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__a21bo_4
MACRO sky130_fd_sc_hd__a21boi_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21boi_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.780000 0.765000 2.170000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.340000 0.765000 2.615000 1.435000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.470000 1.200000 0.895000 1.955000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.392200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.200000 1.610000 1.655000 ;
        RECT 1.065000 1.655000 1.305000 2.465000 ;
        RECT 1.315000 0.255000 1.610000 1.200000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.095000  0.280000 0.380000 0.780000 ;
      RECT 0.095000  0.780000 1.145000 1.030000 ;
      RECT 0.095000  1.030000 0.300000 2.085000 ;
      RECT 0.095000  2.085000 0.355000 2.465000 ;
      RECT 0.525000  2.175000 0.855000 2.635000 ;
      RECT 0.550000  0.085000 1.145000 0.610000 ;
      RECT 1.475000  1.825000 2.665000 2.005000 ;
      RECT 1.475000  2.005000 1.805000 2.465000 ;
      RECT 1.975000  2.175000 2.165000 2.635000 ;
      RECT 2.335000  0.085000 2.665000 0.595000 ;
      RECT 2.335000  2.005000 2.665000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__a21boi_0
MACRO sky130_fd_sc_hd__a21boi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21boi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.760000 0.995000 2.155000 1.345000 ;
        RECT 1.945000 0.375000 2.155000 0.995000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.350000 0.995000 2.640000 1.345000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.975000 0.335000 1.665000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.551000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.045000 1.580000 1.345000 ;
        RECT 1.045000 1.345000 1.375000 2.455000 ;
        RECT 1.335000 0.265000 1.765000 0.795000 ;
        RECT 1.335000 0.795000 1.580000 1.045000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.095000  1.845000 0.855000 2.045000 ;
      RECT 0.095000  2.045000 0.355000 2.435000 ;
      RECT 0.365000  0.265000 0.745000 0.715000 ;
      RECT 0.515000  0.715000 0.745000 1.165000 ;
      RECT 0.515000  1.165000 0.855000 1.845000 ;
      RECT 0.525000  2.225000 0.855000 2.635000 ;
      RECT 0.925000  0.085000 1.155000 0.865000 ;
      RECT 1.545000  1.525000 2.585000 1.725000 ;
      RECT 1.545000  1.725000 1.735000 2.455000 ;
      RECT 1.905000  1.905000 2.235000 2.635000 ;
      RECT 2.325000  0.085000 2.655000 0.815000 ;
      RECT 2.415000  1.725000 2.585000 2.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__a21boi_1
MACRO sky130_fd_sc_hd__a21boi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21boi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.605000 0.995000 3.215000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095000 1.075000 2.425000 1.245000 ;
        RECT 2.100000 1.245000 2.425000 1.495000 ;
        RECT 2.100000 1.495000 3.675000 1.675000 ;
        RECT 3.385000 1.035000 3.795000 1.295000 ;
        RECT 3.385000 1.295000 3.675000 1.495000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.765000 0.425000 1.805000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.627500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.520000 0.255000 1.720000 0.615000 ;
        RECT 1.520000 0.615000 3.060000 0.785000 ;
        RECT 1.520000 0.785000 1.715000 2.115000 ;
        RECT 2.730000 0.255000 3.060000 0.615000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.095000  2.080000 0.425000 2.635000 ;
      RECT 0.265000  0.360000 0.795000 0.530000 ;
      RECT 0.595000  0.530000 0.795000 1.070000 ;
      RECT 0.595000  1.070000 1.325000 1.285000 ;
      RECT 0.595000  1.285000 0.855000 2.265000 ;
      RECT 0.985000  0.085000 1.225000 0.885000 ;
      RECT 1.045000  1.795000 1.350000 2.285000 ;
      RECT 1.045000  2.285000 2.215000 2.465000 ;
      RECT 1.885000  1.855000 3.920000 2.025000 ;
      RECT 1.885000  2.025000 2.215000 2.285000 ;
      RECT 1.940000  0.085000 2.270000 0.445000 ;
      RECT 2.385000  2.195000 2.555000 2.635000 ;
      RECT 2.810000  2.025000 3.920000 2.105000 ;
      RECT 2.810000  2.105000 2.980000 2.465000 ;
      RECT 3.160000  2.275000 3.490000 2.635000 ;
      RECT 3.635000  0.085000 3.930000 0.865000 ;
      RECT 3.660000  2.105000 3.920000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__a21boi_2
MACRO sky130_fd_sc_hd__a21boi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21boi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.545000 1.065000 4.970000 1.310000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.030000 1.065000 3.375000 1.480000 ;
        RECT 3.030000 1.480000 6.450000 1.705000 ;
        RECT 5.205000 1.075000 6.450000 1.480000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 1.075000 0.650000 1.615000 ;
        RECT 0.480000 0.995000 0.650000 1.075000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.288000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.275000 0.370000 1.465000 0.615000 ;
        RECT 1.275000 0.615000 2.325000 0.695000 ;
        RECT 1.275000 0.695000 4.885000 0.865000 ;
        RECT 1.560000 1.585000 2.860000 1.705000 ;
        RECT 1.560000 1.705000 2.725000 2.035000 ;
        RECT 2.135000 0.255000 2.325000 0.615000 ;
        RECT 2.570000 0.865000 4.885000 0.895000 ;
        RECT 2.570000 0.895000 2.860000 1.585000 ;
        RECT 3.255000 0.675000 4.885000 0.695000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.090000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.090000  0.255000 0.445000 0.615000 ;
      RECT 0.090000  0.615000 1.105000 0.795000 ;
      RECT 0.125000  1.785000 0.990000 2.005000 ;
      RECT 0.125000  2.005000 0.455000 2.465000 ;
      RECT 0.625000  2.175000 0.885000 2.635000 ;
      RECT 0.720000  0.085000 1.105000 0.445000 ;
      RECT 0.820000  0.795000 1.105000 1.035000 ;
      RECT 0.820000  1.035000 2.400000 1.345000 ;
      RECT 0.820000  1.345000 0.990000 1.785000 ;
      RECT 1.160000  1.795000 1.355000 2.215000 ;
      RECT 1.160000  2.215000 3.095000 2.465000 ;
      RECT 1.635000  0.085000 1.965000 0.445000 ;
      RECT 1.935000  2.205000 3.095000 2.215000 ;
      RECT 2.495000  0.085000 3.085000 0.525000 ;
      RECT 2.895000  1.875000 6.605000 2.105000 ;
      RECT 2.895000  2.105000 3.095000 2.205000 ;
      RECT 3.265000  0.255000 5.315000 0.505000 ;
      RECT 3.265000  2.275000 3.595000 2.635000 ;
      RECT 4.125000  2.275000 4.455000 2.635000 ;
      RECT 4.625000  2.105000 4.815000 2.465000 ;
      RECT 4.985000  2.275000 5.315000 2.635000 ;
      RECT 5.055000  0.505000 5.315000 0.735000 ;
      RECT 5.055000  0.735000 6.175000 0.905000 ;
      RECT 5.485000  0.085000 5.675000 0.565000 ;
      RECT 5.485000  2.105000 5.665000 2.465000 ;
      RECT 5.845000  0.255000 6.175000 0.735000 ;
      RECT 5.845000  2.275000 6.175000 2.635000 ;
      RECT 6.345000  0.085000 6.605000 0.885000 ;
      RECT 6.345000  2.105000 6.605000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
END sky130_fd_sc_hd__a21boi_4
MACRO sky130_fd_sc_hd__a21o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.660000 1.015000 2.185000 1.325000 ;
        RECT 1.955000 0.375000 2.185000 1.015000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.365000 0.995000 2.665000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 1.015000 1.480000 1.325000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.265000 0.355000 2.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.525000  1.905000 0.865000 2.635000 ;
      RECT 0.545000  0.635000 1.775000 0.835000 ;
      RECT 0.545000  0.835000 0.835000 1.505000 ;
      RECT 0.545000  1.505000 1.315000 1.725000 ;
      RECT 0.615000  0.085000 1.285000 0.455000 ;
      RECT 1.045000  1.725000 1.315000 2.455000 ;
      RECT 1.465000  0.265000 1.775000 0.635000 ;
      RECT 1.495000  1.505000 2.655000 1.745000 ;
      RECT 1.495000  1.745000 1.725000 2.455000 ;
      RECT 1.895000  1.925000 2.225000 2.635000 ;
      RECT 2.365000  0.085000 2.655000 0.815000 ;
      RECT 2.395000  1.745000 2.655000 2.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__a21o_1
MACRO sky130_fd_sc_hd__a21o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.240000 0.365000 2.620000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.810000 0.750000 3.125000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 0.995000 1.790000 1.410000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 0.635000 0.955000 0.825000 ;
        RECT 0.555000 0.825000 0.785000 2.465000 ;
        RECT 0.765000 0.255000 0.955000 0.635000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.095000  1.665000 0.385000 2.635000 ;
      RECT 0.265000  0.085000 0.595000 0.465000 ;
      RECT 0.955000  0.995000 1.295000 1.690000 ;
      RECT 0.955000  1.690000 1.790000 1.920000 ;
      RECT 0.955000  2.220000 1.285000 2.635000 ;
      RECT 1.125000  0.085000 1.455000 0.445000 ;
      RECT 1.125000  0.655000 1.865000 0.825000 ;
      RECT 1.125000  0.825000 1.295000 0.995000 ;
      RECT 1.475000  1.920000 1.790000 2.465000 ;
      RECT 1.675000  0.255000 1.865000 0.655000 ;
      RECT 1.960000  1.670000 3.075000 1.935000 ;
      RECT 1.960000  1.935000 2.185000 2.465000 ;
      RECT 2.355000  2.125000 2.685000 2.635000 ;
      RECT 2.805000  0.085000 3.135000 0.565000 ;
      RECT 2.855000  1.935000 3.075000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a21o_2
MACRO sky130_fd_sc_hd__a21o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.990000 1.010000 4.515000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.425000 1.010000 3.820000 1.275000 ;
        RECT 3.645000 1.275000 3.820000 1.510000 ;
        RECT 3.645000 1.510000 4.935000 1.680000 ;
        RECT 4.685000 1.055000 5.100000 1.290000 ;
        RECT 4.685000 1.290000 4.935000 1.510000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.395000 0.995000 2.705000 1.525000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.615000 1.735000 0.785000 ;
        RECT 0.145000 0.785000 0.630000 1.585000 ;
        RECT 0.145000 1.585000 1.735000 1.755000 ;
        RECT 0.625000 1.755000 0.795000 2.185000 ;
        RECT 1.485000 1.755000 1.735000 2.185000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.105000  0.085000 0.445000 0.445000 ;
      RECT 0.115000  1.935000 0.445000 2.635000 ;
      RECT 0.800000  0.995000 2.205000 1.325000 ;
      RECT 0.975000  0.085000 1.305000 0.445000 ;
      RECT 0.975000  1.935000 1.305000 2.635000 ;
      RECT 1.910000  0.085000 2.685000 0.445000 ;
      RECT 1.915000  1.515000 2.165000 2.635000 ;
      RECT 2.035000  0.615000 3.045000 0.670000 ;
      RECT 2.035000  0.670000 4.365000 0.785000 ;
      RECT 2.035000  0.785000 2.205000 0.995000 ;
      RECT 2.455000  1.695000 2.625000 2.295000 ;
      RECT 2.455000  2.295000 3.465000 2.465000 ;
      RECT 2.875000  0.255000 3.045000 0.615000 ;
      RECT 2.875000  0.785000 4.365000 0.840000 ;
      RECT 2.875000  0.840000 3.045000 2.125000 ;
      RECT 3.255000  0.085000 3.585000 0.445000 ;
      RECT 3.285000  1.445000 3.465000 1.850000 ;
      RECT 3.285000  1.850000 5.360000 2.020000 ;
      RECT 3.285000  2.020000 3.465000 2.295000 ;
      RECT 3.635000  2.275000 3.965000 2.635000 ;
      RECT 4.085000  0.405000 4.365000 0.670000 ;
      RECT 4.135000  2.020000 4.305000 2.465000 ;
      RECT 4.475000  2.275000 4.805000 2.635000 ;
      RECT 4.945000  0.085000 5.225000 0.885000 ;
      RECT 5.030000  2.020000 5.360000 2.395000 ;
      RECT 5.105000  1.460000 5.360000 1.850000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__a21o_4
MACRO sky130_fd_sc_hd__a21oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.850000 0.995000 1.265000 1.325000 ;
        RECT 1.035000 0.375000 1.265000 0.995000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445000 0.995000 1.740000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.675000 0.335000 1.325000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.447000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.495000 0.680000 1.685000 ;
        RECT 0.095000 1.685000 0.370000 2.455000 ;
        RECT 0.505000 0.645000 0.835000 0.825000 ;
        RECT 0.505000 0.825000 0.680000 1.495000 ;
        RECT 0.610000 0.265000 0.835000 0.645000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.110000  0.085000 0.440000 0.475000 ;
      RECT 0.540000  1.855000 1.745000 2.025000 ;
      RECT 0.540000  2.025000 0.870000 2.455000 ;
      RECT 0.850000  1.525000 1.745000 1.855000 ;
      RECT 1.040000  2.195000 1.235000 2.635000 ;
      RECT 1.415000  2.025000 1.745000 2.455000 ;
      RECT 1.445000  0.085000 1.745000 0.815000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__a21oi_1
MACRO sky130_fd_sc_hd__a21oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.815000 0.995000 1.425000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 1.035000 0.645000 1.495000 ;
        RECT 0.145000 1.495000 1.930000 1.675000 ;
        RECT 1.605000 1.075000 1.935000 1.245000 ;
        RECT 1.605000 1.245000 1.930000 1.495000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.800000 0.995000 3.075000 1.625000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.627500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 0.255000 1.300000 0.615000 ;
        RECT 0.955000 0.615000 2.615000 0.785000 ;
        RECT 2.295000 0.255000 2.615000 0.615000 ;
        RECT 2.315000 0.785000 2.615000 2.115000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.100000  0.085000 0.395000 0.865000 ;
      RECT 0.110000  1.855000 2.145000 2.025000 ;
      RECT 0.110000  2.025000 1.220000 2.105000 ;
      RECT 0.110000  2.105000 0.370000 2.465000 ;
      RECT 0.540000  2.275000 0.870000 2.635000 ;
      RECT 1.050000  2.105000 1.220000 2.465000 ;
      RECT 1.475000  2.195000 1.645000 2.635000 ;
      RECT 1.760000  0.085000 2.090000 0.445000 ;
      RECT 1.815000  2.025000 2.145000 2.285000 ;
      RECT 1.815000  2.285000 3.090000 2.465000 ;
      RECT 2.785000  1.795000 3.090000 2.285000 ;
      RECT 2.795000  0.085000 3.125000 0.825000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a21oi_2
MACRO sky130_fd_sc_hd__a21oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.565000 1.065000 4.000000 1.310000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.050000 1.065000 2.395000 1.480000 ;
        RECT 2.050000 1.480000 5.470000 1.705000 ;
        RECT 4.225000 1.075000 5.470000 1.480000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.400000 1.035000 ;
        RECT 0.090000 1.035000 1.430000 1.415000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.288000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.580000 1.585000 1.880000 1.705000 ;
        RECT 0.580000 1.705000 1.745000 2.035000 ;
        RECT 0.595000 0.370000 0.785000 0.615000 ;
        RECT 0.595000 0.615000 1.645000 0.695000 ;
        RECT 0.595000 0.695000 3.905000 0.865000 ;
        RECT 1.455000 0.255000 1.645000 0.615000 ;
        RECT 1.600000 0.865000 3.905000 0.895000 ;
        RECT 1.600000 0.895000 1.880000 1.585000 ;
        RECT 2.275000 0.675000 3.905000 0.695000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.805000 ;
      RECT 0.180000  1.795000 0.375000 2.215000 ;
      RECT 0.180000  2.215000 2.115000 2.465000 ;
      RECT 0.955000  0.085000 1.285000 0.445000 ;
      RECT 0.955000  2.205000 2.115000 2.215000 ;
      RECT 1.835000  0.085000 2.115000 0.525000 ;
      RECT 1.915000  1.875000 5.625000 2.105000 ;
      RECT 1.915000  2.105000 2.115000 2.205000 ;
      RECT 2.285000  0.255000 4.335000 0.505000 ;
      RECT 2.285000  2.275000 2.615000 2.635000 ;
      RECT 2.785000  2.105000 2.975000 2.465000 ;
      RECT 3.145000  2.275000 3.475000 2.635000 ;
      RECT 3.645000  2.105000 3.835000 2.465000 ;
      RECT 4.005000  2.275000 4.335000 2.635000 ;
      RECT 4.075000  0.505000 4.335000 0.735000 ;
      RECT 4.075000  0.735000 5.195000 0.905000 ;
      RECT 4.505000  0.085000 4.695000 0.565000 ;
      RECT 4.505000  2.105000 4.685000 2.465000 ;
      RECT 4.865000  0.255000 5.195000 0.735000 ;
      RECT 4.865000  2.275000 5.195000 2.635000 ;
      RECT 5.365000  0.085000 5.625000 0.885000 ;
      RECT 5.365000  2.105000 5.625000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__a21oi_4
MACRO sky130_fd_sc_hd__a22o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 0.675000 1.695000 1.075000 ;
        RECT 1.485000 1.075000 1.815000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 1.040000 2.395000 1.345000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.765000 1.075000 1.240000 1.285000 ;
        RECT 1.020000 0.675000 1.240000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.575000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875000 0.255000 3.135000 0.585000 ;
        RECT 2.875000 1.785000 3.135000 2.465000 ;
        RECT 2.965000 0.585000 3.135000 1.785000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  0.085000 0.545000 0.850000 ;
      RECT 0.090000  1.455000 1.265000 1.515000 ;
      RECT 0.090000  1.515000 2.795000 1.625000 ;
      RECT 0.090000  1.625000 0.345000 2.245000 ;
      RECT 0.090000  2.245000 0.425000 2.465000 ;
      RECT 0.595000  1.795000 0.780000 1.885000 ;
      RECT 0.595000  1.885000 2.205000 2.085000 ;
      RECT 0.595000  2.085000 0.825000 2.125000 ;
      RECT 0.820000  0.255000 2.120000 0.465000 ;
      RECT 0.935000  1.625000 2.735000 1.685000 ;
      RECT 0.935000  1.685000 1.265000 1.715000 ;
      RECT 1.370000  1.875000 2.205000 1.885000 ;
      RECT 1.430000  2.255000 1.785000 2.635000 ;
      RECT 1.950000  0.465000 2.120000 0.615000 ;
      RECT 1.950000  0.615000 2.705000 0.740000 ;
      RECT 1.950000  0.740000 2.795000 0.785000 ;
      RECT 1.955000  2.085000 2.205000 2.465000 ;
      RECT 2.375000  0.085000 2.705000 0.445000 ;
      RECT 2.455000  1.855000 2.705000 2.635000 ;
      RECT 2.525000  0.785000 2.795000 0.905000 ;
      RECT 2.595000  1.480000 2.795000 1.515000 ;
      RECT 2.625000  0.905000 2.795000 1.480000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a22o_1
MACRO sky130_fd_sc_hd__a22o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.510000 0.675000 1.720000 1.075000 ;
        RECT 1.510000 1.075000 1.840000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.010000 1.075000 2.415000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.765000 1.075000 1.240000 1.285000 ;
        RECT 1.020000 0.675000 1.240000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.575000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.900000 0.255000 3.160000 0.585000 ;
        RECT 2.900000 1.785000 3.160000 2.465000 ;
        RECT 2.990000 0.585000 3.160000 1.785000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.095000  0.085000 0.545000 0.850000 ;
      RECT 0.095000  1.455000 2.815000 1.625000 ;
      RECT 0.095000  1.625000 0.425000 2.295000 ;
      RECT 0.095000  2.295000 1.265000 2.465000 ;
      RECT 0.595000  1.795000 2.230000 2.035000 ;
      RECT 0.595000  2.035000 0.825000 2.125000 ;
      RECT 0.820000  0.255000 2.145000 0.505000 ;
      RECT 0.935000  2.255000 1.265000 2.295000 ;
      RECT 1.455000  2.215000 1.810000 2.635000 ;
      RECT 1.975000  0.505000 2.145000 0.735000 ;
      RECT 1.975000  0.735000 2.815000 0.905000 ;
      RECT 1.980000  2.035000 2.230000 2.465000 ;
      RECT 2.355000  0.085000 2.685000 0.565000 ;
      RECT 2.400000  1.875000 2.730000 2.635000 ;
      RECT 2.645000  0.905000 2.815000 1.455000 ;
      RECT 3.330000  0.085000 3.500000 0.985000 ;
      RECT 3.330000  1.445000 3.500000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a22o_2
MACRO sky130_fd_sc_hd__a22o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.900000 1.075000 5.395000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.350000 1.075000 4.680000 1.445000 ;
        RECT 4.350000 1.445000 5.735000 1.615000 ;
        RECT 5.565000 1.075000 6.355000 1.275000 ;
        RECT 5.565000 1.275000 5.735000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.125000 1.075000 3.680000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.420000 1.075000 2.955000 1.445000 ;
        RECT 2.420000 1.445000 4.180000 1.615000 ;
        RECT 3.850000 1.075000 4.180000 1.445000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.725000 1.770000 0.905000 ;
        RECT 0.085000 0.905000 0.370000 1.445000 ;
        RECT 0.085000 1.445000 1.730000 1.615000 ;
        RECT 0.600000 0.265000 0.930000 0.725000 ;
        RECT 0.640000 1.615000 0.890000 2.465000 ;
        RECT 1.440000 0.255000 1.770000 0.725000 ;
        RECT 1.480000 1.615000 1.730000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.220000  1.825000 0.470000 2.635000 ;
      RECT 0.260000  0.085000 0.430000 0.555000 ;
      RECT 0.540000  1.075000 2.230000 1.275000 ;
      RECT 1.060000  1.795000 1.310000 2.635000 ;
      RECT 1.100000  0.085000 1.270000 0.555000 ;
      RECT 1.900000  1.275000 2.230000 1.785000 ;
      RECT 1.900000  1.785000 3.930000 1.955000 ;
      RECT 1.900000  2.125000 2.150000 2.635000 ;
      RECT 1.940000  0.085000 2.630000 0.555000 ;
      RECT 1.940000  0.735000 5.310000 0.905000 ;
      RECT 1.940000  0.905000 2.230000 1.075000 ;
      RECT 2.420000  2.125000 2.670000 2.295000 ;
      RECT 2.420000  2.295000 4.430000 2.465000 ;
      RECT 2.800000  0.255000 3.970000 0.475000 ;
      RECT 2.840000  1.955000 3.090000 2.125000 ;
      RECT 3.170000  0.645000 3.605000 0.735000 ;
      RECT 3.260000  2.125000 3.510000 2.295000 ;
      RECT 3.680000  1.955000 3.930000 2.125000 ;
      RECT 4.100000  1.785000 6.110000 1.955000 ;
      RECT 4.100000  1.955000 4.430000 2.295000 ;
      RECT 4.185000  0.085000 4.355000 0.555000 ;
      RECT 4.560000  0.255000 5.730000 0.475000 ;
      RECT 4.600000  2.125000 4.850000 2.635000 ;
      RECT 4.935000  0.645000 5.310000 0.735000 ;
      RECT 5.020000  1.955000 5.270000 2.465000 ;
      RECT 5.440000  2.125000 5.690000 2.635000 ;
      RECT 5.480000  0.475000 5.730000 0.895000 ;
      RECT 5.900000  0.085000 6.070000 0.895000 ;
      RECT 5.905000  1.455000 6.110000 1.785000 ;
      RECT 5.905000  1.955000 6.110000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__a22o_4
MACRO sky130_fd_sc_hd__a22oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.490000 0.675000 1.700000 1.075000 ;
        RECT 1.490000 1.075000 1.840000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.010000 0.995000 2.335000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.765000 1.075000 1.240000 1.275000 ;
        RECT 0.990000 0.675000 1.240000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.765000 0.575000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.858000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.445000 1.840000 1.495000 ;
        RECT 0.095000 1.495000 2.675000 1.625000 ;
        RECT 0.095000 1.625000 0.425000 2.295000 ;
        RECT 0.095000 2.295000 1.265000 2.465000 ;
        RECT 0.820000 0.255000 2.125000 0.505000 ;
        RECT 0.935000 2.255000 1.265000 2.295000 ;
        RECT 1.615000 1.625000 2.675000 1.665000 ;
        RECT 1.945000 0.505000 2.125000 0.655000 ;
        RECT 1.945000 0.655000 2.675000 0.825000 ;
        RECT 2.505000 0.825000 2.675000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.095000  0.085000 0.545000 0.595000 ;
      RECT 0.595000  1.795000 1.475000 1.835000 ;
      RECT 0.595000  1.835000 2.125000 2.035000 ;
      RECT 0.595000  2.035000 1.210000 2.085000 ;
      RECT 0.595000  2.085000 0.825000 2.125000 ;
      RECT 1.435000  2.255000 1.810000 2.635000 ;
      RECT 1.955000  2.035000 2.125000 2.165000 ;
      RECT 2.305000  0.085000 2.635000 0.485000 ;
      RECT 2.360000  1.855000 2.625000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__a22oi_1
MACRO sky130_fd_sc_hd__a22oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.075000 3.100000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.390000 1.075000 4.500000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 1.075000 1.700000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 1.075000 0.780000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.141000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.485000 2.160000 1.655000 ;
        RECT 0.095000 1.655000 0.345000 2.465000 ;
        RECT 0.935000 1.655000 1.265000 2.125000 ;
        RECT 1.355000 0.675000 3.045000 0.845000 ;
        RECT 1.775000 1.655000 2.160000 2.125000 ;
        RECT 1.870000 0.845000 2.160000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.095000  0.255000 0.345000 0.680000 ;
      RECT 0.095000  0.680000 1.185000 0.850000 ;
      RECT 0.515000  0.085000 0.845000 0.510000 ;
      RECT 0.515000  1.825000 0.765000 2.295000 ;
      RECT 0.515000  2.295000 2.625000 2.465000 ;
      RECT 1.015000  0.255000 2.105000 0.505000 ;
      RECT 1.015000  0.505000 1.185000 0.680000 ;
      RECT 1.435000  1.825000 1.605000 2.295000 ;
      RECT 2.295000  0.255000 3.385000 0.505000 ;
      RECT 2.375000  1.485000 4.305000 1.655000 ;
      RECT 2.375000  1.655000 2.625000 2.295000 ;
      RECT 2.795000  1.825000 2.965000 2.635000 ;
      RECT 3.135000  1.655000 3.465000 2.465000 ;
      RECT 3.215000  0.505000 3.385000 0.680000 ;
      RECT 3.215000  0.680000 4.375000 0.850000 ;
      RECT 3.555000  0.085000 3.885000 0.510000 ;
      RECT 3.635000  1.825000 3.805000 2.635000 ;
      RECT 3.975000  1.655000 4.305000 2.465000 ;
      RECT 4.055000  0.255000 4.375000 0.680000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__a22oi_2
MACRO sky130_fd_sc_hd__a22oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.275000 1.075000 5.685000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.910000 1.075000 7.735000 1.285000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615000 1.075000 4.040000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.895000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 1.445000 3.325000 1.625000 ;
        RECT 0.595000 1.625000 0.805000 2.125000 ;
        RECT 1.395000 1.625000 1.645000 2.125000 ;
        RECT 2.195000 0.645000 5.565000 0.885000 ;
        RECT 2.195000 0.885000 2.445000 1.445000 ;
        RECT 2.235000 1.625000 2.485000 2.125000 ;
        RECT 3.075000 1.625000 3.325000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.090000  1.455000 0.425000 2.295000 ;
      RECT 0.090000  2.295000 4.265000 2.465000 ;
      RECT 0.095000  0.255000 0.425000 0.725000 ;
      RECT 0.095000  0.725000 2.025000 0.905000 ;
      RECT 0.595000  0.085000 0.765000 0.555000 ;
      RECT 0.935000  0.255000 1.265000 0.725000 ;
      RECT 0.975000  1.795000 1.225000 2.295000 ;
      RECT 1.435000  0.085000 1.605000 0.555000 ;
      RECT 1.775000  0.255000 3.785000 0.475000 ;
      RECT 1.775000  0.475000 2.025000 0.725000 ;
      RECT 1.815000  1.795000 2.065000 2.295000 ;
      RECT 2.655000  1.795000 2.905000 2.295000 ;
      RECT 3.495000  1.455000 7.625000 1.625000 ;
      RECT 3.495000  1.625000 4.265000 2.295000 ;
      RECT 3.975000  0.255000 5.985000 0.475000 ;
      RECT 4.435000  1.795000 4.685000 2.635000 ;
      RECT 4.855000  1.625000 5.105000 2.465000 ;
      RECT 5.275000  1.795000 5.525000 2.635000 ;
      RECT 5.695000  1.625000 5.945000 2.465000 ;
      RECT 5.735000  0.475000 5.985000 0.725000 ;
      RECT 5.735000  0.725000 7.665000 0.905000 ;
      RECT 6.115000  1.795000 6.365000 2.635000 ;
      RECT 6.155000  0.085000 6.325000 0.555000 ;
      RECT 6.495000  0.255000 6.825000 0.725000 ;
      RECT 6.535000  1.625000 6.785000 2.465000 ;
      RECT 6.955000  1.795000 7.205000 2.635000 ;
      RECT 6.995000  0.085000 7.165000 0.555000 ;
      RECT 7.335000  0.255000 7.665000 0.725000 ;
      RECT 7.375000  1.625000 7.625000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__a22oi_4
MACRO sky130_fd_sc_hd__a31o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895000 0.995000 2.160000 1.655000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 0.995000 1.700000 1.655000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935000 0.995000 1.240000 1.325000 ;
        RECT 1.025000 1.325000 1.240000 1.655000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 0.995000 2.620000 1.655000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.437250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.300000 0.425000 0.810000 ;
        RECT 0.095000 0.810000 0.285000 1.575000 ;
        RECT 0.095000 1.575000 0.425000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.455000  0.995000 0.765000 1.325000 ;
      RECT 0.595000  0.085000 0.925000 0.485000 ;
      RECT 0.595000  0.655000 2.960000 0.825000 ;
      RECT 0.595000  0.825000 0.765000 0.995000 ;
      RECT 0.595000  1.495000 0.845000 2.635000 ;
      RECT 1.035000  1.825000 2.325000 1.995000 ;
      RECT 1.035000  1.995000 1.285000 2.415000 ;
      RECT 1.515000  2.165000 1.845000 2.635000 ;
      RECT 1.975000  0.315000 2.305000 0.655000 ;
      RECT 2.075000  1.995000 2.325000 2.415000 ;
      RECT 2.475000  0.085000 2.805000 0.485000 ;
      RECT 2.505000  1.825000 2.960000 1.995000 ;
      RECT 2.505000  1.995000 2.835000 2.425000 ;
      RECT 2.790000  0.825000 2.960000 1.825000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a31o_1
MACRO sky130_fd_sc_hd__a31o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 0.415000 2.175000 0.700000 ;
        RECT 1.965000 0.700000 2.355000 0.870000 ;
        RECT 2.185000 0.870000 2.355000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 0.400000 1.700000 0.695000 ;
        RECT 1.530000 0.695000 1.795000 0.865000 ;
        RECT 1.625000 0.865000 1.795000 1.075000 ;
        RECT 1.625000 1.075000 1.955000 1.245000 ;
        RECT 1.625000 1.245000 1.795000 1.260000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.760000 1.270000 0.995000 ;
        RECT 1.065000 0.995000 1.395000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895000 0.755000 3.090000 1.325000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.715000 0.765000 0.885000 ;
        RECT 0.090000 0.885000 0.345000 1.835000 ;
        RECT 0.090000 1.835000 0.765000 2.005000 ;
        RECT 0.595000 0.255000 0.765000 0.715000 ;
        RECT 0.595000 2.005000 0.765000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  0.085000 0.345000 0.545000 ;
      RECT 0.135000  2.175000 0.385000 2.635000 ;
      RECT 0.555000  1.075000 0.885000 1.245000 ;
      RECT 0.555000  1.245000 0.725000 1.495000 ;
      RECT 0.555000  1.495000 3.045000 1.665000 ;
      RECT 0.935000  1.835000 1.185000 2.635000 ;
      RECT 0.955000  0.085000 1.285000 0.465000 ;
      RECT 1.015000  0.465000 1.185000 0.545000 ;
      RECT 1.355000  1.835000 2.645000 2.005000 ;
      RECT 1.355000  2.005000 1.605000 2.425000 ;
      RECT 1.815000  2.175000 2.145000 2.635000 ;
      RECT 2.335000  2.005000 2.585000 2.425000 ;
      RECT 2.375000  0.335000 2.705000 0.505000 ;
      RECT 2.460000  0.255000 2.705000 0.335000 ;
      RECT 2.535000  0.505000 2.705000 1.495000 ;
      RECT 2.875000  0.085000 3.135000 0.565000 ;
      RECT 2.875000  1.665000 3.045000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a31o_2
MACRO sky130_fd_sc_hd__a31o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.075000 1.705000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.725000 1.075000 1.055000 1.245000 ;
        RECT 0.805000 0.735000 2.170000 0.905000 ;
        RECT 0.805000 0.905000 0.975000 1.075000 ;
        RECT 1.985000 0.905000 2.170000 1.075000 ;
        RECT 1.985000 1.075000 2.315000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 1.075000 0.525000 1.445000 ;
        RECT 0.150000 1.445000 2.855000 1.615000 ;
        RECT 2.525000 1.075000 2.855000 1.445000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.575000 1.075000 4.030000 1.285000 ;
        RECT 3.815000 0.745000 4.030000 1.075000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.505000 0.655000 6.295000 0.825000 ;
        RECT 4.535000 1.785000 6.295000 1.955000 ;
        RECT 4.595000 1.955000 4.765000 2.465000 ;
        RECT 5.435000 1.955000 5.605000 2.465000 ;
        RECT 6.125000 0.825000 6.295000 1.785000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.175000  0.085000 0.345000 0.905000 ;
      RECT 0.175000  1.785000 2.985000 1.955000 ;
      RECT 0.175000  1.955000 0.345000 2.465000 ;
      RECT 0.515000  2.125000 0.845000 2.635000 ;
      RECT 1.015000  1.955000 1.185000 2.465000 ;
      RECT 1.355000  0.395000 2.520000 0.565000 ;
      RECT 1.355000  2.125000 1.685000 2.635000 ;
      RECT 1.855000  1.955000 2.025000 2.465000 ;
      RECT 2.195000  2.125000 2.525000 2.635000 ;
      RECT 2.350000  0.565000 2.520000 0.700000 ;
      RECT 2.350000  0.700000 3.485000 0.805000 ;
      RECT 2.350000  0.805000 3.345000 0.870000 ;
      RECT 2.700000  0.085000 2.985000 0.530000 ;
      RECT 2.815000  1.955000 2.985000 2.295000 ;
      RECT 2.815000  2.295000 3.825000 2.465000 ;
      RECT 3.155000  0.295000 3.485000 0.700000 ;
      RECT 3.155000  0.870000 3.345000 1.455000 ;
      RECT 3.155000  1.455000 4.395000 1.625000 ;
      RECT 3.155000  1.625000 3.485000 2.115000 ;
      RECT 3.655000  1.795000 3.825000 2.295000 ;
      RECT 3.735000  0.085000 4.265000 0.565000 ;
      RECT 4.095000  2.125000 4.425000 2.635000 ;
      RECT 4.225000  0.995000 5.935000 1.325000 ;
      RECT 4.225000  1.325000 4.395000 1.455000 ;
      RECT 4.935000  0.085000 5.265000 0.485000 ;
      RECT 4.935000  2.125000 5.265000 2.635000 ;
      RECT 5.775000  0.085000 6.105000 0.485000 ;
      RECT 5.775000  2.125000 6.105000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__a31o_4
MACRO sky130_fd_sc_hd__a31oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 1.445000 1.455000 1.665000 ;
        RECT 1.270000 0.995000 1.455000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 0.335000 1.055000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.365000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 0.995000 2.215000 1.325000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.481250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.380000 0.295000 1.785000 0.715000 ;
        RECT 1.380000 0.715000 1.795000 0.825000 ;
        RECT 1.625000 0.825000 1.795000 1.495000 ;
        RECT 1.625000 1.495000 2.210000 1.665000 ;
        RECT 1.875000 1.665000 2.210000 2.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.090000  0.085000 0.430000 0.815000 ;
      RECT 0.090000  1.495000 0.420000 2.635000 ;
      RECT 0.590000  1.835000 1.695000 2.005000 ;
      RECT 0.590000  2.005000 0.765000 2.415000 ;
      RECT 0.935000  2.175000 1.265000 2.635000 ;
      RECT 1.470000  2.005000 1.695000 2.415000 ;
      RECT 1.955000  0.085000 2.215000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__a31oi_1
MACRO sky130_fd_sc_hd__a31oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 0.995000 2.665000 1.615000 ;
        RECT 2.905000 0.995000 3.075000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.995000 1.755000 1.615000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.995000 0.820000 1.615000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.820000 1.075000 4.490000 1.275000 ;
        RECT 4.265000 1.275000 4.490000 1.625000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.922000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295000 0.655000 4.505000 0.825000 ;
        RECT 3.255000 0.255000 3.425000 0.655000 ;
        RECT 3.255000 0.825000 3.570000 1.445000 ;
        RECT 3.255000 1.445000 4.085000 1.615000 ;
        RECT 3.755000 1.615000 4.085000 2.115000 ;
        RECT 4.175000 0.295000 4.505000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.095000  0.655000 2.105000 0.825000 ;
      RECT 0.175000  1.785000 3.505000 1.955000 ;
      RECT 0.175000  1.955000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.125000 0.845000 2.635000 ;
      RECT 1.015000  1.955000 1.185000 2.465000 ;
      RECT 1.355000  0.295000 3.075000 0.465000 ;
      RECT 1.355000  2.125000 1.685000 2.635000 ;
      RECT 1.855000  1.955000 2.025000 2.465000 ;
      RECT 2.310000  2.125000 2.980000 2.635000 ;
      RECT 3.335000  1.955000 3.505000 2.295000 ;
      RECT 3.335000  2.295000 4.425000 2.465000 ;
      RECT 3.675000  0.085000 4.005000 0.465000 ;
      RECT 4.255000  1.795000 4.425000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__a31oi_2
MACRO sky130_fd_sc_hd__a31oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825000 0.995000 5.420000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.995000 3.550000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.995000 1.735000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.670000 0.995000 6.855000 1.630000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.443500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.975000 0.635000 7.585000 0.805000 ;
        RECT 6.075000 1.915000 7.245000 2.085000 ;
        RECT 6.575000 0.255000 6.745000 0.635000 ;
        RECT 7.045000 0.805000 7.245000 1.915000 ;
        RECT 7.415000 0.255000 7.585000 0.635000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.175000  0.255000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 3.785000 0.805000 ;
      RECT 0.175000  1.495000 5.405000 1.665000 ;
      RECT 0.175000  1.665000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  1.915000 0.845000 2.635000 ;
      RECT 1.015000  0.255000 1.185000 0.635000 ;
      RECT 1.015000  1.665000 1.185000 2.465000 ;
      RECT 1.355000  0.085000 1.685000 0.465000 ;
      RECT 1.355000  1.915000 1.685000 2.635000 ;
      RECT 1.855000  0.255000 2.025000 0.635000 ;
      RECT 1.855000  1.665000 2.025000 2.465000 ;
      RECT 2.195000  0.295000 5.565000 0.465000 ;
      RECT 2.195000  1.915000 2.525000 2.635000 ;
      RECT 2.695000  1.665000 2.865000 2.465000 ;
      RECT 3.035000  1.915000 3.365000 2.635000 ;
      RECT 3.535000  1.665000 3.705000 2.465000 ;
      RECT 3.895000  1.915000 4.225000 2.635000 ;
      RECT 4.395000  1.665000 4.565000 2.465000 ;
      RECT 4.735000  2.255000 5.065000 2.635000 ;
      RECT 5.235000  1.665000 5.405000 2.255000 ;
      RECT 5.235000  2.255000 7.665000 2.425000 ;
      RECT 5.235000  2.425000 5.405000 2.465000 ;
      RECT 6.075000  0.085000 6.405000 0.465000 ;
      RECT 6.915000  0.085000 7.245000 0.465000 ;
      RECT 7.415000  1.495000 7.665000 2.255000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__a31oi_4
MACRO sky130_fd_sc_hd__a32o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 0.665000 2.280000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 0.665000 1.800000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 0.995000 1.320000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.450000 0.660000 2.870000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.180000 0.995000 3.530000 1.325000 ;
        RECT 3.325000 1.325000 3.530000 1.615000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.544500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.300000 0.425000 0.560000 ;
        RECT 0.090000 0.560000 0.345000 1.915000 ;
        RECT 0.090000 1.915000 0.425000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.570000  0.995000 0.875000 1.325000 ;
      RECT 0.595000  0.085000 0.925000 0.485000 ;
      RECT 0.675000  1.835000 1.005000 2.635000 ;
      RECT 0.705000  0.655000 1.265000 0.825000 ;
      RECT 0.705000  0.825000 0.875000 0.995000 ;
      RECT 0.705000  1.325000 0.875000 1.495000 ;
      RECT 0.705000  1.495000 3.075000 1.665000 ;
      RECT 1.095000  0.315000 2.710000 0.485000 ;
      RECT 1.095000  0.485000 1.265000 0.655000 ;
      RECT 1.250000  1.875000 2.675000 2.045000 ;
      RECT 1.250000  2.045000 1.535000 2.465000 ;
      RECT 1.790000  2.215000 2.120000 2.635000 ;
      RECT 2.345000  2.045000 2.675000 2.295000 ;
      RECT 2.345000  2.295000 3.505000 2.465000 ;
      RECT 2.905000  1.665000 3.075000 2.125000 ;
      RECT 3.255000  0.085000 3.585000 0.805000 ;
      RECT 3.335000  1.795000 3.505000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a32o_1
MACRO sky130_fd_sc_hd__a32o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.685000 0.955000 2.985000 1.325000 ;
        RECT 2.755000 0.415000 3.105000 0.610000 ;
        RECT 2.755000 0.610000 2.985000 0.955000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.165000 0.995000 3.545000 1.325000 ;
        RECT 3.305000 0.425000 3.545000 0.995000 ;
        RECT 3.305000 1.325000 3.545000 1.625000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 0.995000 4.055000 1.630000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.085000 1.075000 2.515000 1.245000 ;
        RECT 2.345000 1.245000 2.515000 1.445000 ;
        RECT 2.345000 1.445000 2.550000 1.615000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 0.745000 1.530000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.695500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 0.655000 0.845000 0.825000 ;
        RECT 0.135000 0.825000 0.345000 1.785000 ;
        RECT 0.135000 1.785000 1.185000 1.955000 ;
        RECT 0.135000 1.955000 0.345000 2.465000 ;
        RECT 1.015000 1.955000 1.185000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.465000 ;
      RECT 0.515000  2.125000 0.845000 2.635000 ;
      RECT 0.535000  0.995000 0.705000 1.445000 ;
      RECT 0.535000  1.445000 2.125000 1.615000 ;
      RECT 0.935000  0.085000 1.640000 0.445000 ;
      RECT 1.535000  1.785000 1.705000 2.295000 ;
      RECT 1.535000  2.295000 2.545000 2.465000 ;
      RECT 1.700000  0.615000 2.585000 0.785000 ;
      RECT 1.700000  0.785000 1.890000 1.445000 ;
      RECT 1.875000  1.615000 2.125000 1.945000 ;
      RECT 1.875000  1.945000 2.205000 2.115000 ;
      RECT 2.255000  0.275000 2.585000 0.615000 ;
      RECT 2.375000  1.795000 3.545000 1.965000 ;
      RECT 2.375000  1.965000 2.545000 2.295000 ;
      RECT 2.715000  2.140000 3.045000 2.635000 ;
      RECT 3.375000  1.965000 3.545000 2.465000 ;
      RECT 3.715000  0.085000 4.050000 0.805000 ;
      RECT 3.715000  1.915000 4.050000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__a32o_2
MACRO sky130_fd_sc_hd__a32o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.280000 1.075000 5.075000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.335000 1.075000 4.030000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.210000 1.075000 3.105000 1.295000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.630000 1.075000 6.780000 1.625000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.030000 1.075000 7.710000 1.295000 ;
        RECT 7.030000 1.295000 7.225000 1.635000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.635000 1.605000 0.805000 ;
        RECT 0.120000 0.805000 0.340000 1.495000 ;
        RECT 0.120000 1.495000 1.605000 1.665000 ;
        RECT 0.595000 0.255000 0.765000 0.635000 ;
        RECT 0.595000 1.665000 0.765000 2.465000 ;
        RECT 1.435000 0.255000 1.605000 0.635000 ;
        RECT 1.435000 1.665000 1.605000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.095000  1.915000 0.425000 2.635000 ;
      RECT 0.570000  0.995000 1.970000 1.325000 ;
      RECT 0.935000  0.085000 1.265000 0.465000 ;
      RECT 0.935000  1.915000 1.265000 2.635000 ;
      RECT 1.775000  0.085000 2.105000 0.465000 ;
      RECT 1.775000  1.915000 2.105000 2.635000 ;
      RECT 1.800000  1.325000 1.970000 1.495000 ;
      RECT 1.800000  1.495000 5.450000 1.665000 ;
      RECT 2.275000  0.255000 2.445000 0.655000 ;
      RECT 2.275000  0.655000 3.885000 0.825000 ;
      RECT 2.275000  1.915000 5.065000 2.085000 ;
      RECT 2.275000  2.085000 2.445000 2.465000 ;
      RECT 2.615000  0.085000 2.945000 0.465000 ;
      RECT 2.615000  2.255000 2.945000 2.635000 ;
      RECT 3.135000  0.295000 5.145000 0.465000 ;
      RECT 3.215000  2.085000 3.385000 2.465000 ;
      RECT 3.555000  2.255000 3.885000 2.635000 ;
      RECT 4.055000  2.085000 4.225000 2.465000 ;
      RECT 4.395000  0.635000 6.425000 0.805000 ;
      RECT 4.395000  2.255000 4.725000 2.635000 ;
      RECT 4.895000  2.085000 5.065000 2.255000 ;
      RECT 4.895000  2.255000 7.725000 2.425000 ;
      RECT 5.280000  0.805000 5.450000 1.495000 ;
      RECT 5.280000  1.665000 5.450000 1.905000 ;
      RECT 5.280000  1.905000 6.200000 1.915000 ;
      RECT 5.280000  1.915000 7.305000 2.075000 ;
      RECT 5.670000  0.295000 6.805000 0.465000 ;
      RECT 6.135000  2.075000 7.305000 2.085000 ;
      RECT 6.635000  0.255000 6.805000 0.295000 ;
      RECT 6.635000  0.465000 6.805000 0.645000 ;
      RECT 6.635000  0.645000 7.645000 0.815000 ;
      RECT 6.975000  0.085000 7.305000 0.465000 ;
      RECT 7.475000  0.255000 7.645000 0.645000 ;
      RECT 7.475000  1.755000 7.725000 2.255000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__a32o_4
MACRO sky130_fd_sc_hd__a32oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.230000 1.075000 1.595000 1.255000 ;
        RECT 1.405000 0.345000 1.705000 0.765000 ;
        RECT 1.405000 0.765000 1.595000 1.075000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 0.995000 2.165000 1.325000 ;
        RECT 1.965000 0.415000 2.165000 0.995000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335000 1.015000 2.750000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 0.995000 1.025000 1.425000 ;
        RECT 0.855000 1.425000 1.255000 1.615000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.345000 1.325000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.575500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.635000 1.165000 0.805000 ;
        RECT 0.515000 0.805000 0.685000 1.785000 ;
        RECT 0.515000 1.785000 0.865000 2.085000 ;
        RECT 0.915000 0.295000 1.165000 0.635000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  1.835000 0.345000 2.255000 ;
      RECT 0.085000  2.255000 1.345000 2.465000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 1.095000  1.785000 2.185000 1.955000 ;
      RECT 1.095000  1.955000 1.345000 2.255000 ;
      RECT 1.555000  2.135000 1.805000 2.635000 ;
      RECT 2.015000  1.745000 2.185000 1.785000 ;
      RECT 2.015000  1.955000 2.185000 2.465000 ;
      RECT 2.355000  0.085000 2.695000 0.805000 ;
      RECT 2.355000  1.495000 2.695000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a32oi_1
MACRO sky130_fd_sc_hd__a32oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415000 1.075000 3.220000 1.625000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725000 1.075000 4.480000 1.625000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.715000 1.075000 5.860000 1.625000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.080000 1.725000 1.285000 ;
        RECT 1.175000 1.075000 1.505000 1.080000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 1.075000 0.825000 1.285000 ;
        RECT 0.145000 1.285000 0.325000 1.625000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.955000 0.845000 2.125000 ;
        RECT 0.595000 1.455000 2.180000 1.625000 ;
        RECT 0.595000 1.625000 0.765000 1.955000 ;
        RECT 1.355000 0.655000 3.100000 0.825000 ;
        RECT 1.435000 1.625000 1.605000 2.125000 ;
        RECT 1.965000 0.825000 2.180000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.095000  0.295000 0.425000 0.465000 ;
      RECT 0.175000  0.465000 0.345000 0.715000 ;
      RECT 0.175000  0.715000 1.185000 0.885000 ;
      RECT 0.175000  1.795000 0.345000 2.295000 ;
      RECT 0.175000  2.295000 2.025000 2.465000 ;
      RECT 0.595000  0.085000 0.765000 0.545000 ;
      RECT 0.935000  0.295000 2.115000 0.465000 ;
      RECT 1.015000  0.465000 1.185000 0.715000 ;
      RECT 1.015000  1.795000 1.185000 2.295000 ;
      RECT 1.855000  1.795000 2.025000 1.915000 ;
      RECT 1.855000  1.915000 5.805000 2.085000 ;
      RECT 1.855000  2.085000 2.025000 2.295000 ;
      RECT 2.270000  2.255000 2.940000 2.635000 ;
      RECT 2.350000  0.295000 4.370000 0.465000 ;
      RECT 3.180000  1.795000 3.350000 1.915000 ;
      RECT 3.180000  2.085000 3.350000 2.465000 ;
      RECT 3.550000  2.255000 4.220000 2.635000 ;
      RECT 3.620000  0.635000 5.390000 0.805000 ;
      RECT 4.390000  1.795000 4.560000 1.915000 ;
      RECT 4.390000  2.085000 4.560000 2.465000 ;
      RECT 4.555000  0.085000 4.890000 0.465000 ;
      RECT 4.765000  2.255000 5.435000 2.635000 ;
      RECT 5.060000  0.275000 5.390000 0.635000 ;
      RECT 5.560000  0.085000 5.885000 0.885000 ;
      RECT 5.635000  1.795000 5.805000 1.915000 ;
      RECT 5.635000  2.085000 5.805000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__a32oi_2
MACRO sky130_fd_sc_hd__a32oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775000 1.075000 5.465000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.095000 1.075000 7.695000 1.300000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.295000 1.075000 9.985000 1.280000 ;
        RECT 9.805000 0.755000 9.985000 1.075000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.585000 0.995000 3.555000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 1.750000 1.305000 ;
        RECT 0.110000 1.305000 0.330000 1.965000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.575000 3.365000 1.745000 ;
        RECT 0.515000 1.745000 0.845000 2.085000 ;
        RECT 1.355000 1.745000 1.685000 2.085000 ;
        RECT 1.975000 0.990000 2.365000 1.575000 ;
        RECT 1.975000 1.745000 2.525000 2.085000 ;
        RECT 2.195000 0.635000 5.565000 0.805000 ;
        RECT 2.195000 0.805000 2.365000 0.990000 ;
        RECT 3.035000 1.745000 3.365000 2.085000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.095000  2.255000  3.705000 2.425000 ;
      RECT 0.175000  0.255000  0.345000 0.635000 ;
      RECT 0.175000  0.635000  2.025000 0.805000 ;
      RECT 0.515000  0.085000  0.845000 0.465000 ;
      RECT 1.015000  0.255000  1.185000 0.635000 ;
      RECT 1.355000  0.085000  1.685000 0.465000 ;
      RECT 1.855000  0.295000  3.785000 0.465000 ;
      RECT 1.855000  0.465000  2.025000 0.635000 ;
      RECT 3.535000  1.575000  9.925000 1.745000 ;
      RECT 3.535000  1.745000  3.705000 2.255000 ;
      RECT 3.895000  1.915000  4.225000 2.635000 ;
      RECT 3.975000  0.295000  7.805000 0.465000 ;
      RECT 4.395000  1.745000  4.565000 2.465000 ;
      RECT 4.770000  1.915000  5.440000 2.635000 ;
      RECT 5.640000  1.745000  5.810000 2.465000 ;
      RECT 6.215000  0.635000  9.505000 0.805000 ;
      RECT 6.215000  1.915000  6.545000 2.635000 ;
      RECT 6.715000  1.745000  6.885000 2.465000 ;
      RECT 7.055000  1.915000  7.385000 2.635000 ;
      RECT 7.555000  1.745000  7.725000 2.465000 ;
      RECT 7.995000  0.085000  8.325000 0.465000 ;
      RECT 8.415000  1.915000  8.745000 2.635000 ;
      RECT 8.495000  0.255000  8.665000 0.635000 ;
      RECT 8.835000  0.085000  9.165000 0.465000 ;
      RECT 8.915000  1.745000  9.085000 2.465000 ;
      RECT 9.255000  1.915000  9.585000 2.635000 ;
      RECT 9.335000  0.255000  9.505000 0.635000 ;
      RECT 9.685000  0.085000 10.025000 0.465000 ;
      RECT 9.755000  1.745000  9.925000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
END sky130_fd_sc_hd__a32oi_4
MACRO sky130_fd_sc_hd__a41o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 0.995000 1.915000 1.325000 ;
        RECT 1.535000 1.325000 1.835000 1.620000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.700000 0.415000 2.650000 0.600000 ;
        RECT 2.225000 0.600000 2.445000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.705000 0.995000 3.085000 1.625000 ;
        RECT 2.880000 0.395000 3.085000 0.995000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 0.995000 3.570000 1.625000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.075000 1.335000 1.635000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.300000 0.425000 0.560000 ;
        RECT 0.085000 0.560000 0.345000 2.165000 ;
        RECT 0.085000 2.165000 0.425000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.515000  0.735000 1.530000 0.810000 ;
      RECT 0.515000  0.810000 1.335000 0.905000 ;
      RECT 0.515000  0.905000 0.685000 1.825000 ;
      RECT 0.515000  1.825000 1.365000 1.995000 ;
      RECT 0.595000  0.085000 0.925000 0.565000 ;
      RECT 0.595000  2.175000 0.845000 2.635000 ;
      RECT 1.035000  1.995000 1.365000 2.425000 ;
      RECT 1.115000  0.300000 1.530000 0.735000 ;
      RECT 1.535000  1.795000 3.505000 1.965000 ;
      RECT 1.535000  1.965000 1.705000 2.465000 ;
      RECT 1.915000  2.175000 2.165000 2.635000 ;
      RECT 2.375000  1.965000 2.545000 2.465000 ;
      RECT 2.845000  2.175000 3.095000 2.635000 ;
      RECT 3.255000  0.085000 3.595000 0.810000 ;
      RECT 3.335000  1.965000 3.505000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a41o_1
MACRO sky130_fd_sc_hd__a41o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.785000 0.730000 4.005000 1.625000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.085000 1.075000 3.550000 1.245000 ;
        RECT 3.335000 0.745000 3.550000 1.075000 ;
        RECT 3.335000 1.245000 3.550000 1.625000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.685000 0.995000 2.855000 1.435000 ;
        RECT 2.685000 1.435000 3.090000 1.625000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.000000 0.995000 2.335000 1.625000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.400000 1.075000 1.730000 1.295000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.295000 0.765000 0.755000 ;
        RECT 0.595000 0.755000 0.785000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.805000 ;
      RECT 0.095000  1.495000 0.425000 2.635000 ;
      RECT 0.935000  0.085000 1.265000 0.465000 ;
      RECT 0.980000  0.635000 2.545000 0.805000 ;
      RECT 0.980000  0.805000 1.150000 1.495000 ;
      RECT 0.980000  1.495000 1.785000 1.665000 ;
      RECT 1.015000  1.835000 1.265000 2.635000 ;
      RECT 1.455000  1.665000 1.785000 2.425000 ;
      RECT 1.495000  0.255000 1.705000 0.635000 ;
      RECT 1.875000  0.085000 2.205000 0.465000 ;
      RECT 1.955000  1.795000 3.965000 1.965000 ;
      RECT 1.955000  1.965000 2.125000 2.465000 ;
      RECT 2.335000  2.175000 2.585000 2.635000 ;
      RECT 2.375000  0.295000 4.045000 0.465000 ;
      RECT 2.375000  0.465000 2.545000 0.635000 ;
      RECT 2.795000  1.965000 2.965000 2.465000 ;
      RECT 3.335000  2.175000 3.585000 2.635000 ;
      RECT 3.795000  1.965000 3.965000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__a41o_2
MACRO sky130_fd_sc_hd__a41o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395000 1.075000 4.065000 1.295000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.275000 1.075000 4.975000 1.285000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.155000 1.075000 6.185000 1.295000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.495000 1.075000 7.505000 1.295000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.135000 1.075000 3.145000 1.280000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.635000 1.605000 0.805000 ;
        RECT 0.150000 0.805000 0.320000 1.575000 ;
        RECT 0.150000 1.575000 1.605000 1.745000 ;
        RECT 0.595000 0.255000 0.765000 0.635000 ;
        RECT 0.595000 1.745000 0.765000 2.465000 ;
        RECT 1.435000 0.255000 1.605000 0.635000 ;
        RECT 1.435000 1.745000 1.605000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.095000  1.915000 0.425000 2.635000 ;
      RECT 0.490000  1.075000 1.945000 1.245000 ;
      RECT 0.935000  0.085000 1.265000 0.465000 ;
      RECT 0.935000  1.915000 1.265000 2.635000 ;
      RECT 1.775000  0.085000 2.125000 0.465000 ;
      RECT 1.775000  0.645000 3.905000 0.815000 ;
      RECT 1.775000  0.815000 1.945000 1.075000 ;
      RECT 1.775000  1.245000 1.945000 1.455000 ;
      RECT 1.775000  1.455000 2.965000 1.625000 ;
      RECT 1.775000  1.915000 2.125000 2.635000 ;
      RECT 2.295000  0.255000 2.465000 0.645000 ;
      RECT 2.375000  1.795000 2.545000 2.295000 ;
      RECT 2.375000  2.295000 3.405000 2.465000 ;
      RECT 2.635000  0.085000 2.965000 0.465000 ;
      RECT 2.715000  1.955000 3.045000 2.125000 ;
      RECT 2.795000  1.625000 2.965000 1.955000 ;
      RECT 3.155000  0.295000 4.245000 0.465000 ;
      RECT 3.235000  1.535000 7.370000 1.705000 ;
      RECT 3.235000  1.705000 3.405000 2.295000 ;
      RECT 3.575000  1.915000 3.905000 2.635000 ;
      RECT 4.075000  0.465000 4.245000 0.645000 ;
      RECT 4.075000  0.645000 5.165000 0.815000 ;
      RECT 4.075000  1.705000 4.245000 2.465000 ;
      RECT 4.415000  0.295000 6.105000 0.465000 ;
      RECT 4.415000  1.915000 4.745000 2.635000 ;
      RECT 4.935000  1.705000 5.105000 2.465000 ;
      RECT 5.345000  1.915000 6.035000 2.635000 ;
      RECT 5.355000  0.645000 7.285000 0.815000 ;
      RECT 6.275000  1.705000 6.445000 2.465000 ;
      RECT 6.615000  0.085000 6.945000 0.465000 ;
      RECT 6.615000  1.915000 6.945000 2.635000 ;
      RECT 7.115000  0.255000 7.285000 0.645000 ;
      RECT 7.115000  1.705000 7.285000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__a41o_4
MACRO sky130_fd_sc_hd__a41oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.780000 0.995000 3.085000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.890000 0.755000 2.210000 1.665000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.470000 0.755000 1.710000 1.665000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.960000 0.965000 1.250000 1.665000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 0.965000 0.780000 1.665000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.669500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.285000 0.345000 0.615000 ;
        RECT 0.090000 0.615000 1.290000 0.785000 ;
        RECT 0.090000 0.785000 0.360000 1.845000 ;
        RECT 0.090000 1.845000 0.425000 2.425000 ;
        RECT 1.120000 0.295000 3.015000 0.465000 ;
        RECT 1.120000 0.465000 1.290000 0.615000 ;
        RECT 2.685000 0.465000 3.015000 0.805000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.595000  1.845000 3.015000 2.015000 ;
      RECT 0.595000  2.015000 0.845000 2.465000 ;
      RECT 0.620000  0.085000 0.950000 0.445000 ;
      RECT 1.120000  2.195000 1.450000 2.635000 ;
      RECT 1.760000  2.015000 1.930000 2.465000 ;
      RECT 2.215000  2.195000 2.545000 2.635000 ;
      RECT 2.765000  2.015000 3.015000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a41oi_1
MACRO sky130_fd_sc_hd__a41oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.785000 1.075000 2.455000 1.295000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.665000 1.075000 3.365000 1.285000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.545000 1.075000 4.575000 1.295000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.755000 1.075000 5.895000 1.295000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.075000 1.555000 1.280000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.645000 2.295000 0.815000 ;
        RECT 0.145000 0.815000 0.315000 1.455000 ;
        RECT 0.145000 1.455000 1.455000 1.625000 ;
        RECT 0.685000 0.255000 0.855000 0.645000 ;
        RECT 1.125000 1.625000 1.455000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.185000  0.085000 0.515000 0.465000 ;
      RECT 0.785000  1.795000 0.955000 2.295000 ;
      RECT 0.785000  2.295000 1.795000 2.465000 ;
      RECT 1.025000  0.085000 1.375000 0.465000 ;
      RECT 1.545000  0.295000 2.635000 0.465000 ;
      RECT 1.625000  1.535000 5.760000 1.705000 ;
      RECT 1.625000  1.705000 1.795000 2.295000 ;
      RECT 1.965000  1.915000 2.295000 2.635000 ;
      RECT 2.465000  0.465000 2.635000 0.645000 ;
      RECT 2.465000  0.645000 3.555000 0.815000 ;
      RECT 2.465000  1.705000 2.635000 2.465000 ;
      RECT 2.805000  0.295000 4.495000 0.465000 ;
      RECT 2.805000  1.915000 3.135000 2.635000 ;
      RECT 3.325000  1.705000 3.495000 2.465000 ;
      RECT 3.745000  0.645000 5.675000 0.815000 ;
      RECT 3.755000  1.915000 4.425000 2.635000 ;
      RECT 4.665000  1.705000 4.835000 2.465000 ;
      RECT 5.005000  0.085000 5.335000 0.465000 ;
      RECT 5.005000  1.915000 5.335000 2.635000 ;
      RECT 5.505000  0.255000 5.675000 0.645000 ;
      RECT 5.505000  1.705000 5.675000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__a41oi_2
MACRO sky130_fd_sc_hd__a41oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.385000 0.995000 4.205000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.405000 1.075000 6.315000 1.285000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.560000 1.075000 7.955000 1.300000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285000 1.075000 9.975000 1.280000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 1.745000 1.305000 ;
        RECT 0.105000 1.305000 0.325000 1.965000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.575000 2.155000 1.685000 ;
        RECT 0.515000 1.685000 1.685000 1.745000 ;
        RECT 0.515000 1.745000 0.845000 2.085000 ;
        RECT 0.595000 0.255000 0.765000 0.635000 ;
        RECT 0.595000 0.635000 4.015000 0.805000 ;
        RECT 1.350000 1.495000 2.155000 1.575000 ;
        RECT 1.350000 1.745000 1.685000 2.085000 ;
        RECT 1.435000 0.255000 1.605000 0.635000 ;
        RECT 1.935000 0.805000 2.155000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.090000  0.085000  0.425000 0.465000 ;
      RECT 0.090000  2.255000  2.335000 2.425000 ;
      RECT 0.935000  0.085000  1.265000 0.465000 ;
      RECT 1.775000  0.085000  2.105000 0.465000 ;
      RECT 2.165000  1.905000  3.515000 2.075000 ;
      RECT 2.165000  2.075000  2.335000 2.255000 ;
      RECT 2.165000  2.425000  2.335000 2.465000 ;
      RECT 2.425000  0.295000  6.115000 0.465000 ;
      RECT 2.505000  2.255000  3.175000 2.635000 ;
      RECT 3.345000  1.575000  9.945000 1.745000 ;
      RECT 3.345000  1.745000  3.515000 1.905000 ;
      RECT 3.345000  2.075000  3.515000 2.465000 ;
      RECT 3.685000  1.915000  4.015000 2.635000 ;
      RECT 4.185000  1.745000  4.355000 2.425000 ;
      RECT 4.525000  0.635000  7.895000 0.805000 ;
      RECT 4.620000  1.915000  4.950000 2.635000 ;
      RECT 5.120000  1.745000  5.290000 2.465000 ;
      RECT 5.495000  1.915000  6.165000 2.635000 ;
      RECT 6.305000  0.295000  8.235000 0.465000 ;
      RECT 6.385000  1.745000  6.555000 2.465000 ;
      RECT 6.725000  1.915000  7.055000 2.635000 ;
      RECT 7.225000  1.745000  7.395000 2.465000 ;
      RECT 7.565000  1.915000  7.895000 2.635000 ;
      RECT 8.065000  0.255000  8.235000 0.295000 ;
      RECT 8.065000  0.465000  8.235000 0.635000 ;
      RECT 8.065000  0.635000  9.915000 0.805000 ;
      RECT 8.065000  1.745000  8.235000 2.465000 ;
      RECT 8.405000  0.085000  8.735000 0.465000 ;
      RECT 8.405000  1.915000  8.735000 2.635000 ;
      RECT 8.905000  0.255000  9.075000 0.635000 ;
      RECT 8.905000  1.745000  9.075000 2.465000 ;
      RECT 9.245000  0.085000  9.575000 0.465000 ;
      RECT 9.245000  1.915000  9.575000 2.635000 ;
      RECT 9.745000  0.255000  9.915000 0.635000 ;
      RECT 9.775000  1.745000  9.945000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
END sky130_fd_sc_hd__a41oi_4
MACRO sky130_fd_sc_hd__a211o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 0.995000 2.060000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 0.995000 1.305000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.240000 0.995000 2.675000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855000 0.995000 3.125000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.437250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.265000 0.425000 1.685000 ;
        RECT 0.090000 1.685000 0.355000 2.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.135000 -0.085000 0.305000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.525000  1.915000 0.855000 2.635000 ;
      RECT 0.600000  0.625000 3.085000 0.815000 ;
      RECT 0.600000  0.815000 0.825000 1.505000 ;
      RECT 0.600000  1.505000 3.095000 1.685000 ;
      RECT 0.605000  0.085000 1.350000 0.455000 ;
      RECT 1.045000  1.865000 2.235000 2.095000 ;
      RECT 1.045000  2.095000 1.305000 2.455000 ;
      RECT 1.475000  2.265000 1.805000 2.635000 ;
      RECT 1.915000  0.265000 2.170000 0.625000 ;
      RECT 1.975000  2.095000 2.235000 2.455000 ;
      RECT 2.350000  0.085000 2.680000 0.455000 ;
      RECT 2.805000  1.685000 3.095000 2.455000 ;
      RECT 2.860000  0.265000 3.085000 0.625000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a211o_1
MACRO sky130_fd_sc_hd__a211o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.980000 1.045000 2.450000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 1.045000 1.810000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.620000 1.045000 3.070000 1.275000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.260000 1.045000 3.595000 1.275000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.452000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 0.255000 0.775000 0.635000 ;
        RECT 0.555000 0.635000 0.785000 2.335000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.090000  0.085000 0.385000 0.905000 ;
      RECT 0.090000  1.490000 0.385000 2.635000 ;
      RECT 0.945000  0.085000 1.795000 0.445000 ;
      RECT 1.000000  0.695000 3.585000 0.875000 ;
      RECT 1.000000  0.875000 1.310000 1.490000 ;
      RECT 1.000000  1.490000 3.585000 1.660000 ;
      RECT 1.000000  1.830000 1.255000 2.635000 ;
      RECT 1.455000  1.840000 2.795000 2.020000 ;
      RECT 1.455000  2.020000 1.785000 2.465000 ;
      RECT 1.955000  2.190000 2.230000 2.635000 ;
      RECT 2.275000  0.275000 2.605000 0.695000 ;
      RECT 2.465000  2.020000 2.795000 2.465000 ;
      RECT 2.810000  0.085000 3.085000 0.525000 ;
      RECT 3.255000  0.275000 3.585000 0.695000 ;
      RECT 3.255000  1.660000 3.585000 2.325000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a211o_2
MACRO sky130_fd_sc_hd__a211o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.035000 1.020000 5.380000 1.330000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.495000 1.020000 4.825000 1.510000 ;
        RECT 4.495000 1.510000 5.845000 1.700000 ;
        RECT 5.635000 1.020000 6.225000 1.320000 ;
        RECT 5.635000 1.320000 5.845000 1.510000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.540000 0.985000 2.805000 1.325000 ;
        RECT 2.625000 1.325000 2.805000 1.445000 ;
        RECT 2.625000 1.445000 4.175000 1.700000 ;
        RECT 3.845000 0.985000 4.175000 1.445000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.975000 0.985000 3.645000 1.275000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.933750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.635000 2.025000 0.875000 ;
        RECT 0.085000 0.875000 0.340000 1.495000 ;
        RECT 0.085000 1.495000 1.640000 1.705000 ;
        RECT 0.595000 1.705000 0.780000 2.465000 ;
        RECT 0.985000 0.255000 1.175000 0.615000 ;
        RECT 0.985000 0.615000 2.025000 0.635000 ;
        RECT 1.450000 1.705000 1.640000 2.465000 ;
        RECT 1.845000 0.255000 2.025000 0.615000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.090000  1.875000 0.425000 2.635000 ;
      RECT 0.485000  0.085000 0.815000 0.465000 ;
      RECT 0.525000  1.045000 2.370000 1.325000 ;
      RECT 0.950000  1.875000 1.280000 2.635000 ;
      RECT 1.345000  0.085000 1.675000 0.445000 ;
      RECT 1.810000  1.835000 2.060000 2.635000 ;
      RECT 2.185000  1.325000 2.370000 1.505000 ;
      RECT 2.185000  1.505000 2.455000 1.675000 ;
      RECT 2.195000  0.615000 5.490000 0.805000 ;
      RECT 2.195000  0.805000 2.370000 1.045000 ;
      RECT 2.220000  0.085000 2.555000 0.445000 ;
      RECT 2.280000  1.675000 2.455000 1.870000 ;
      RECT 2.280000  1.870000 3.510000 2.040000 ;
      RECT 2.320000  2.210000 4.450000 2.465000 ;
      RECT 2.725000  0.255000 2.970000 0.615000 ;
      RECT 3.140000  0.085000 3.470000 0.445000 ;
      RECT 3.640000  0.255000 4.020000 0.615000 ;
      RECT 4.120000  1.880000 6.345000 2.105000 ;
      RECT 4.120000  2.105000 4.450000 2.210000 ;
      RECT 4.190000  0.085000 4.560000 0.445000 ;
      RECT 4.620000  2.275000 4.950000 2.635000 ;
      RECT 5.160000  0.275000 5.490000 0.615000 ;
      RECT 5.160000  2.105000 5.420000 2.465000 ;
      RECT 5.590000  2.275000 5.920000 2.635000 ;
      RECT 6.015000  0.085000 6.345000 0.805000 ;
      RECT 6.015000  1.535000 6.345000 1.880000 ;
      RECT 6.090000  2.105000 6.345000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__a211o_4
MACRO sky130_fd_sc_hd__a211oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.265000 0.855000 0.995000 ;
        RECT 0.605000 0.995000 1.245000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.765000 0.435000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.425000 0.995000 1.755000 1.325000 ;
        RECT 1.525000 1.325000 1.755000 2.455000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.995000 2.235000 1.615000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.619250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.180000 0.265000 1.365000 0.625000 ;
        RECT 1.180000 0.625000 2.660000 0.815000 ;
        RECT 1.935000 1.785000 2.660000 2.455000 ;
        RECT 2.055000 0.265000 2.280000 0.625000 ;
        RECT 2.445000 0.815000 2.660000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.085000 0.425000 0.595000 ;
      RECT 0.250000  1.525000 1.355000 1.725000 ;
      RECT 0.250000  1.725000 0.500000 2.455000 ;
      RECT 0.670000  1.905000 1.000000 2.635000 ;
      RECT 1.170000  1.725000 1.355000 2.455000 ;
      RECT 1.545000  0.085000 1.875000 0.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__a211oi_1
MACRO sky130_fd_sc_hd__a211oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.370000 1.035000 3.080000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.740000 1.035000 4.500000 1.285000 ;
        RECT 4.175000 1.285000 4.500000 1.655000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 1.035000 1.785000 1.285000 ;
        RECT 1.035000 1.285000 1.255000 1.615000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.995000 0.405000 1.615000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.826000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575000 0.255000 0.835000 0.655000 ;
        RECT 0.575000 0.655000 3.145000 0.855000 ;
        RECT 0.575000 0.855000 0.855000 1.785000 ;
        RECT 0.575000 1.785000 0.905000 2.105000 ;
        RECT 1.505000 0.285000 1.695000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.125000 -0.085000 0.295000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.145000  0.085000 0.395000 0.815000 ;
      RECT 0.145000  1.785000 0.405000 2.285000 ;
      RECT 0.145000  2.285000 2.215000 2.455000 ;
      RECT 1.005000  0.085000 1.335000 0.475000 ;
      RECT 1.075000  1.785000 1.265000 2.255000 ;
      RECT 1.075000  2.255000 2.215000 2.285000 ;
      RECT 1.435000  1.455000 3.975000 1.655000 ;
      RECT 1.435000  1.655000 1.765000 2.075000 ;
      RECT 1.865000  0.085000 2.195000 0.475000 ;
      RECT 1.935000  1.835000 2.215000 2.255000 ;
      RECT 2.385000  0.265000 3.495000 0.475000 ;
      RECT 2.435000  1.835000 2.665000 2.635000 ;
      RECT 2.845000  1.655000 3.115000 2.465000 ;
      RECT 3.295000  1.835000 3.525000 2.635000 ;
      RECT 3.325000  0.475000 3.495000 0.635000 ;
      RECT 3.325000  0.635000 4.435000 0.855000 ;
      RECT 3.675000  0.085000 4.005000 0.455000 ;
      RECT 3.705000  1.655000 3.975000 2.465000 ;
      RECT 4.155000  1.835000 4.385000 2.635000 ;
      RECT 4.185000  0.265000 4.435000 0.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__a211oi_2
MACRO sky130_fd_sc_hd__a211oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655000 1.075000 3.005000 1.245000 ;
        RECT 1.660000 1.035000 3.005000 1.075000 ;
        RECT 1.660000 1.245000 3.005000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.035000 1.385000 1.445000 ;
        RECT 0.100000 1.445000 3.575000 1.625000 ;
        RECT 3.245000 1.035000 3.575000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.745000 1.035000 4.755000 1.275000 ;
        RECT 3.745000 1.275000 4.460000 1.615000 ;
      LAYER mcon ;
        RECT 3.830000 1.445000 4.000000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.590000 0.995000 6.935000 1.325000 ;
        RECT 6.590000 1.325000 6.760000 1.615000 ;
      LAYER mcon ;
        RECT 6.590000 1.445000 6.760000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.770000 1.415000 4.060000 1.460000 ;
        RECT 3.770000 1.460000 6.820000 1.600000 ;
        RECT 3.770000 1.600000 4.060000 1.645000 ;
        RECT 6.530000 1.415000 6.820000 1.460000 ;
        RECT 6.530000 1.600000 6.820000 1.645000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.000000 1.035000 6.350000 1.275000 ;
        RECT 6.130000 1.275000 6.350000 1.695000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.685000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775000 0.675000 3.330000 0.695000 ;
        RECT 1.775000 0.695000 7.275000 0.825000 ;
        RECT 1.775000 0.825000 6.355000 0.865000 ;
        RECT 3.875000 0.255000 4.195000 0.615000 ;
        RECT 3.875000 0.615000 5.045000 0.625000 ;
        RECT 3.875000 0.625000 7.275000 0.695000 ;
        RECT 4.875000 0.255000 5.045000 0.615000 ;
        RECT 5.170000 1.865000 7.275000 2.085000 ;
        RECT 5.715000 0.255000 5.885000 0.615000 ;
        RECT 5.715000 0.615000 7.275000 0.625000 ;
        RECT 6.930000 1.495000 7.275000 1.865000 ;
        RECT 7.105000 0.825000 7.275000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.095000  0.085000 0.395000 0.585000 ;
      RECT 0.095000  1.795000 3.705000 2.085000 ;
      RECT 0.095000  2.085000 0.345000 2.465000 ;
      RECT 0.515000  2.255000 0.845000 2.635000 ;
      RECT 0.565000  0.530000 0.775000 0.695000 ;
      RECT 0.565000  0.695000 1.605000 0.865000 ;
      RECT 0.950000  0.085000 1.185000 0.525000 ;
      RECT 1.015000  2.085000 3.705000 2.105000 ;
      RECT 1.015000  2.105000 1.185000 2.465000 ;
      RECT 1.355000  0.255000 3.365000 0.505000 ;
      RECT 1.355000  0.505000 1.605000 0.695000 ;
      RECT 1.355000  2.275000 1.685000 2.635000 ;
      RECT 1.855000  2.105000 2.025000 2.465000 ;
      RECT 2.195000  2.275000 2.525000 2.635000 ;
      RECT 2.695000  2.105000 2.865000 2.465000 ;
      RECT 3.035000  2.275000 3.365000 2.635000 ;
      RECT 3.535000  0.085000 3.705000 0.525000 ;
      RECT 3.535000  2.105000 3.705000 2.255000 ;
      RECT 3.535000  2.255000 7.270000 2.465000 ;
      RECT 3.875000  1.785000 4.910000 2.085000 ;
      RECT 4.365000  0.085000 4.695000 0.445000 ;
      RECT 4.630000  1.445000 5.960000 1.695000 ;
      RECT 4.630000  1.695000 4.910000 1.785000 ;
      RECT 5.215000  0.085000 5.545000 0.445000 ;
      RECT 6.055000  0.085000 6.385000 0.445000 ;
      RECT 6.915000  0.085000 7.270000 0.445000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__a211oi_4
MACRO sky130_fd_sc_hd__a221o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.970000 0.675000 2.255000 1.075000 ;
        RECT 1.970000 1.075000 2.300000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.470000 1.075000 2.835000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225000 1.075000 1.700000 1.275000 ;
        RECT 1.420000 0.675000 1.700000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 1.075000 1.055000 1.275000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.440000 1.285000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.320000 0.255000 3.575000 0.585000 ;
        RECT 3.320000 1.795000 3.575000 2.465000 ;
        RECT 3.390000 0.585000 3.575000 0.665000 ;
        RECT 3.405000 0.665000 3.575000 1.795000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.175000  0.255000 0.345000 0.735000 ;
      RECT 0.175000  0.735000 1.240000 0.905000 ;
      RECT 0.175000  1.455000 3.235000 1.625000 ;
      RECT 0.175000  1.625000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.565000 ;
      RECT 0.515000  1.795000 0.845000 2.295000 ;
      RECT 0.515000  2.295000 1.685000 2.465000 ;
      RECT 1.015000  1.795000 2.650000 2.035000 ;
      RECT 1.015000  2.035000 1.245000 2.125000 ;
      RECT 1.070000  0.255000 2.605000 0.505000 ;
      RECT 1.070000  0.505000 1.240000 0.735000 ;
      RECT 1.355000  2.255000 1.685000 2.295000 ;
      RECT 1.875000  2.215000 2.230000 2.635000 ;
      RECT 2.400000  2.035000 2.650000 2.465000 ;
      RECT 2.435000  0.505000 2.605000 0.735000 ;
      RECT 2.435000  0.735000 3.235000 0.905000 ;
      RECT 2.775000  0.085000 3.105000 0.565000 ;
      RECT 2.820000  1.875000 3.150000 2.635000 ;
      RECT 3.065000  0.905000 3.235000 1.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a221o_1
MACRO sky130_fd_sc_hd__a221o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.970000 0.675000 2.255000 1.075000 ;
        RECT 1.970000 1.075000 2.300000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.470000 1.075000 2.835000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225000 1.075000 1.700000 1.275000 ;
        RECT 1.420000 0.675000 1.700000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 1.075000 1.055000 1.275000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.440000 1.285000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.320000 0.255000 3.575000 0.585000 ;
        RECT 3.320000 1.795000 3.575000 2.465000 ;
        RECT 3.390000 0.585000 3.575000 0.665000 ;
        RECT 3.405000 0.665000 3.575000 1.795000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.175000  0.255000 0.345000 0.735000 ;
      RECT 0.175000  0.735000 1.240000 0.905000 ;
      RECT 0.175000  1.455000 3.235000 1.625000 ;
      RECT 0.175000  1.625000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.565000 ;
      RECT 0.515000  1.795000 0.845000 2.295000 ;
      RECT 0.515000  2.295000 1.685000 2.465000 ;
      RECT 1.015000  1.795000 2.650000 2.035000 ;
      RECT 1.015000  2.035000 1.245000 2.125000 ;
      RECT 1.070000  0.255000 2.605000 0.505000 ;
      RECT 1.070000  0.505000 1.240000 0.735000 ;
      RECT 1.355000  2.255000 1.685000 2.295000 ;
      RECT 1.875000  2.215000 2.230000 2.635000 ;
      RECT 2.400000  2.035000 2.650000 2.465000 ;
      RECT 2.435000  0.505000 2.605000 0.735000 ;
      RECT 2.435000  0.735000 3.235000 0.905000 ;
      RECT 2.775000  0.085000 3.105000 0.565000 ;
      RECT 2.820000  1.875000 3.150000 2.635000 ;
      RECT 3.065000  0.905000 3.235000 1.455000 ;
      RECT 3.745000  0.085000 3.915000 0.980000 ;
      RECT 3.745000  1.445000 3.915000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__a221o_2
MACRO sky130_fd_sc_hd__a221o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855000 1.075000 3.190000 1.105000 ;
        RECT 2.855000 1.105000 4.060000 1.285000 ;
        RECT 3.710000 1.075000 4.060000 1.105000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.265000 1.075000 2.680000 1.285000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235000 1.075000 6.035000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.270000 1.075000 7.280000 1.285000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.230000 1.075000 4.725000 1.285000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.735000 1.685000 0.905000 ;
        RECT 0.095000 0.905000 0.325000 1.455000 ;
        RECT 0.095000 1.455000 1.645000 1.625000 ;
        RECT 0.515000 0.255000 0.845000 0.725000 ;
        RECT 0.515000 0.725000 1.685000 0.735000 ;
        RECT 0.555000 1.625000 0.805000 2.465000 ;
        RECT 1.355000 0.255000 1.685000 0.725000 ;
        RECT 1.395000 1.625000 1.645000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.155000  1.795000 0.385000 2.635000 ;
      RECT 0.175000  0.085000 0.345000 0.555000 ;
      RECT 0.495000  1.075000 1.845000 1.115000 ;
      RECT 0.495000  1.115000 1.985000 1.285000 ;
      RECT 0.975000  1.795000 1.225000 2.635000 ;
      RECT 1.015000  0.085000 1.185000 0.555000 ;
      RECT 1.815000  1.285000 1.985000 1.455000 ;
      RECT 1.815000  1.455000 5.065000 1.625000 ;
      RECT 1.815000  1.795000 2.065000 2.635000 ;
      RECT 1.855000  0.085000 2.025000 0.555000 ;
      RECT 1.855000  0.735000 2.525000 0.905000 ;
      RECT 1.945000  0.905000 2.165000 0.935000 ;
      RECT 2.195000  0.255000 2.525000 0.735000 ;
      RECT 2.235000  1.795000 4.230000 1.875000 ;
      RECT 2.235000  1.875000 5.575000 1.965000 ;
      RECT 2.235000  1.965000 2.485000 2.465000 ;
      RECT 2.655000  2.135000 2.905000 2.635000 ;
      RECT 2.695000  0.085000 2.865000 0.895000 ;
      RECT 3.075000  1.965000 3.330000 2.465000 ;
      RECT 3.080000  0.305000 4.305000 0.475000 ;
      RECT 3.190000  0.735000 3.885000 0.905000 ;
      RECT 3.315000  0.905000 3.610000 0.935000 ;
      RECT 3.500000  2.135000 3.750000 2.635000 ;
      RECT 3.550000  0.645000 3.885000 0.735000 ;
      RECT 3.940000  2.215000 6.385000 2.295000 ;
      RECT 3.940000  2.295000 7.225000 2.465000 ;
      RECT 4.055000  0.475000 4.305000 0.725000 ;
      RECT 4.055000  0.725000 5.065000 0.905000 ;
      RECT 4.060000  1.965000 5.575000 2.045000 ;
      RECT 4.405000  1.625000 4.735000 1.705000 ;
      RECT 4.475000  0.085000 4.645000 0.555000 ;
      RECT 4.815000  0.255000 5.985000 0.475000 ;
      RECT 4.815000  0.475000 5.065000 0.725000 ;
      RECT 4.895000  0.905000 5.065000 1.455000 ;
      RECT 5.235000  0.645000 6.505000 0.725000 ;
      RECT 5.235000  0.725000 7.345000 0.905000 ;
      RECT 5.245000  1.455000 6.805000 1.625000 ;
      RECT 5.245000  1.625000 5.575000 1.875000 ;
      RECT 5.745000  1.795000 6.385000 2.215000 ;
      RECT 6.555000  1.625000 6.805000 2.125000 ;
      RECT 6.675000  0.085000 6.845000 0.555000 ;
      RECT 6.975000  1.785000 7.225000 2.295000 ;
      RECT 7.015000  0.255000 7.345000 0.725000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 1.995000  0.765000 2.165000 0.935000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.400000  0.765000 3.570000 0.935000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 1.935000 0.735000 2.225000 0.780000 ;
      RECT 1.935000 0.780000 3.630000 0.920000 ;
      RECT 1.935000 0.920000 2.225000 0.965000 ;
      RECT 3.340000 0.735000 3.630000 0.780000 ;
      RECT 3.340000 0.920000 3.630000 0.965000 ;
  END
END sky130_fd_sc_hd__a221o_4
MACRO sky130_fd_sc_hd__a221oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 0.675000 2.200000 1.075000 ;
        RECT 1.945000 1.075000 2.275000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.470000 0.995000 2.755000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225000 1.075000 1.695000 1.285000 ;
        RECT 1.415000 0.675000 1.695000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 1.075000 1.055000 1.285000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.435000 1.285000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.767000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.170000 0.255000 0.345000 0.735000 ;
        RECT 0.170000 0.735000 1.235000 0.905000 ;
        RECT 0.175000 1.455000 2.300000 1.495000 ;
        RECT 0.175000 1.495000 3.135000 1.625000 ;
        RECT 0.175000 1.625000 0.345000 2.465000 ;
        RECT 1.065000 0.255000 2.580000 0.505000 ;
        RECT 1.065000 0.505000 1.235000 0.735000 ;
        RECT 2.150000 1.625000 3.135000 1.665000 ;
        RECT 2.380000 0.505000 2.580000 0.655000 ;
        RECT 2.380000 0.655000 3.135000 0.825000 ;
        RECT 2.925000 0.825000 3.135000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.515000  0.085000 0.845000 0.565000 ;
      RECT 0.515000  1.795000 0.765000 2.295000 ;
      RECT 0.515000  2.295000 1.685000 2.465000 ;
      RECT 1.015000  1.795000 2.025000 1.835000 ;
      RECT 1.015000  1.835000 2.625000 2.045000 ;
      RECT 1.015000  2.045000 1.240000 2.125000 ;
      RECT 1.355000  2.255000 1.685000 2.295000 ;
      RECT 1.875000  2.215000 2.205000 2.635000 ;
      RECT 2.375000  2.045000 2.625000 2.465000 ;
      RECT 2.750000  0.085000 3.080000 0.485000 ;
      RECT 2.795000  1.875000 3.125000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a221oi_1
MACRO sky130_fd_sc_hd__a221oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.985000 1.075000 4.480000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.435000 1.075000 3.765000 1.445000 ;
        RECT 3.435000 1.445000 4.820000 1.615000 ;
        RECT 4.650000 1.075000 5.435000 1.275000 ;
        RECT 4.650000 1.275000 4.820000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.210000 1.075000 2.765000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.075000 2.040000 1.445000 ;
        RECT 1.505000 1.445000 3.265000 1.615000 ;
        RECT 2.935000 1.075000 3.265000 1.445000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.420000 1.615000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.796500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 0.305000 0.855000 0.725000 ;
        RECT 0.525000 0.725000 4.395000 0.865000 ;
        RECT 0.605000 0.865000 4.395000 0.905000 ;
        RECT 0.605000 0.905000 0.855000 2.125000 ;
        RECT 2.285000 0.645000 2.635000 0.725000 ;
        RECT 4.065000 0.645000 4.395000 0.725000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.090000  1.795000 0.435000 2.295000 ;
      RECT 0.090000  2.295000 1.275000 2.465000 ;
      RECT 0.105000  0.085000 0.355000 0.895000 ;
      RECT 1.025000  0.085000 1.715000 0.555000 ;
      RECT 1.025000  1.495000 1.275000 1.785000 ;
      RECT 1.025000  1.785000 3.015000 1.955000 ;
      RECT 1.025000  1.955000 1.275000 2.295000 ;
      RECT 1.505000  2.125000 1.755000 2.295000 ;
      RECT 1.505000  2.295000 3.475000 2.465000 ;
      RECT 1.885000  0.255000 3.055000 0.475000 ;
      RECT 1.925000  1.955000 2.175000 2.125000 ;
      RECT 2.345000  2.125000 2.595000 2.295000 ;
      RECT 2.765000  1.955000 3.015000 2.125000 ;
      RECT 3.225000  1.785000 5.195000 1.955000 ;
      RECT 3.225000  1.955000 3.475000 2.295000 ;
      RECT 3.270000  0.085000 3.440000 0.555000 ;
      RECT 3.645000  0.255000 4.815000 0.475000 ;
      RECT 3.685000  2.125000 3.935000 2.635000 ;
      RECT 4.105000  1.955000 4.355000 2.465000 ;
      RECT 4.525000  2.125000 4.775000 2.635000 ;
      RECT 4.565000  0.475000 4.815000 0.905000 ;
      RECT 4.985000  0.085000 5.155000 0.905000 ;
      RECT 4.990000  1.455000 5.195000 1.785000 ;
      RECT 4.990000  1.955000 5.195000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__a221oi_2
MACRO sky130_fd_sc_hd__a221oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.475000 1.075000 7.885000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.965000 1.075000 6.295000 1.445000 ;
        RECT 5.965000 1.445000 8.265000 1.615000 ;
        RECT 8.095000 1.075000 9.575000 1.275000 ;
        RECT 8.095000 1.275000 8.265000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.935000 0.995000 5.285000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.415000 0.995000 3.765000 1.325000 ;
        RECT 3.595000 1.325000 3.765000 1.445000 ;
        RECT 3.595000 1.445000 5.795000 1.615000 ;
        RECT 5.465000 1.075000 5.795000 1.445000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.335000 1.275000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.593000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 1.705000 0.905000 ;
        RECT 0.575000 1.445000 1.705000 1.615000 ;
        RECT 0.575000 1.615000 0.825000 2.125000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 1.415000 1.615000 1.665000 2.125000 ;
        RECT 1.505000 0.905000 1.705000 1.095000 ;
        RECT 1.505000 1.095000 3.245000 1.275000 ;
        RECT 1.505000 1.275000 1.705000 1.445000 ;
        RECT 3.075000 0.645000 5.680000 0.735000 ;
        RECT 3.075000 0.735000 7.765000 0.820000 ;
        RECT 3.075000 0.820000 3.245000 1.095000 ;
        RECT 5.510000 0.820000 6.460000 0.905000 ;
        RECT 6.290000 0.645000 7.765000 0.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.090000  1.445000 0.405000 2.295000 ;
      RECT 0.090000  2.295000 2.125000 2.465000 ;
      RECT 0.115000  0.085000 0.365000 0.895000 ;
      RECT 0.995000  1.785000 1.245000 2.295000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.875000  0.085000 2.045000 0.645000 ;
      RECT 1.875000  0.645000 2.905000 0.925000 ;
      RECT 1.875000  1.445000 3.030000 1.615000 ;
      RECT 1.875000  1.615000 2.125000 2.295000 ;
      RECT 2.235000  0.255000 5.585000 0.425000 ;
      RECT 2.235000  0.425000 2.610000 0.475000 ;
      RECT 2.315000  1.795000 2.565000 2.215000 ;
      RECT 2.315000  2.215000 6.005000 2.465000 ;
      RECT 2.735000  0.595000 2.905000 0.645000 ;
      RECT 2.735000  1.615000 3.030000 1.835000 ;
      RECT 2.735000  1.835000 5.585000 2.045000 ;
      RECT 3.035000  0.425000 5.585000 0.475000 ;
      RECT 5.755000  1.785000 8.605000 2.045000 ;
      RECT 5.755000  2.045000 6.005000 2.215000 ;
      RECT 5.835000  0.085000 6.005000 0.555000 ;
      RECT 6.175000  0.255000 8.185000 0.475000 ;
      RECT 6.175000  2.215000 8.185000 2.635000 ;
      RECT 7.935000  0.475000 8.185000 0.725000 ;
      RECT 7.935000  0.725000 9.025000 0.905000 ;
      RECT 8.355000  0.085000 8.525000 0.555000 ;
      RECT 8.355000  2.045000 8.525000 2.465000 ;
      RECT 8.435000  1.445000 9.405000 1.615000 ;
      RECT 8.435000  1.615000 8.605000 1.785000 ;
      RECT 8.695000  0.255000 9.025000 0.725000 ;
      RECT 8.775000  1.795000 8.945000 2.635000 ;
      RECT 9.155000  1.615000 9.405000 2.465000 ;
      RECT 9.195000  0.085000 9.365000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
END sky130_fd_sc_hd__a221oi_4
MACRO sky130_fd_sc_hd__a222oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a222oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615000 1.000000 2.925000 1.330000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095000 1.000000 3.435000 1.330000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.135000 1.000000 2.445000 1.330000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655000 1.000000 1.965000 1.330000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.000000 0.545000 1.315000 ;
    END
  END C1
  PIN C2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.715000 1.000000 1.085000 1.315000 ;
    END
  END C2
  PIN Y
    ANTENNADIFFAREA  0.897600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.255000 0.425000 0.645000 ;
        RECT 0.095000 0.645000 2.645000 0.815000 ;
        RECT 0.095000 1.485000 0.425000 1.500000 ;
        RECT 0.095000 1.500000 1.425000 1.670000 ;
        RECT 0.095000 1.670000 0.425000 1.680000 ;
        RECT 0.095000 1.680000 0.345000 2.255000 ;
        RECT 0.095000 2.255000 0.425000 2.465000 ;
        RECT 1.015000 1.670000 1.185000 1.830000 ;
        RECT 1.255000 0.815000 1.480000 1.330000 ;
        RECT 1.255000 1.330000 1.425000 1.500000 ;
        RECT 2.315000 0.295000 2.645000 0.645000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 3.680000 0.240000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.515000  1.875000 0.845000 2.075000 ;
      RECT 0.595000  2.075000 0.765000 2.295000 ;
      RECT 0.595000  2.295000 2.185000 2.465000 ;
      RECT 0.875000  0.085000 1.605000 0.465000 ;
      RECT 1.515000  1.825000 2.015000 1.965000 ;
      RECT 1.515000  1.965000 1.970000 1.970000 ;
      RECT 1.515000  1.970000 1.935000 1.980000 ;
      RECT 1.515000  1.980000 1.915000 1.995000 ;
      RECT 1.845000  1.655000 3.595000 1.670000 ;
      RECT 1.845000  1.670000 2.685000 1.735000 ;
      RECT 1.845000  1.735000 2.605000 1.825000 ;
      RECT 2.015000  2.135000 2.185000 2.295000 ;
      RECT 2.355000  1.500000 3.595000 1.655000 ;
      RECT 2.355000  1.825000 2.605000 2.255000 ;
      RECT 2.355000  2.255000 2.685000 2.465000 ;
      RECT 2.775000  1.905000 3.105000 2.075000 ;
      RECT 2.855000  2.075000 3.025000 2.635000 ;
      RECT 3.220000  1.670000 3.595000 1.735000 ;
      RECT 3.255000  0.085000 3.585000 0.815000 ;
      RECT 3.255000  2.255000 3.595000 2.465000 ;
      RECT 3.335000  1.735000 3.595000 2.255000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a222oi_1
MACRO sky130_fd_sc_hd__a311o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 0.765000 2.155000 0.995000 ;
        RECT 1.965000 0.995000 2.310000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.510000 0.750000 1.705000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.905000 0.995000 1.240000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.620000 0.995000 3.095000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.350000 0.995000 3.535000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.454000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.395000 0.670000 ;
        RECT 0.085000 0.670000 0.255000 1.785000 ;
        RECT 0.085000 1.785000 0.425000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.425000  0.995000 0.735000 1.325000 ;
      RECT 0.565000  0.655000 1.260000 0.825000 ;
      RECT 0.565000  0.825000 0.735000 0.995000 ;
      RECT 0.565000  1.325000 0.735000 1.495000 ;
      RECT 0.565000  1.495000 3.505000 1.665000 ;
      RECT 0.590000  0.085000 0.920000 0.465000 ;
      RECT 0.595000  2.175000 0.840000 2.635000 ;
      RECT 1.015000  1.835000 2.575000 2.005000 ;
      RECT 1.015000  2.005000 1.265000 2.465000 ;
      RECT 1.090000  0.255000 2.495000 0.425000 ;
      RECT 1.090000  0.425000 1.260000 0.655000 ;
      RECT 1.455000  2.255000 2.125000 2.635000 ;
      RECT 2.325000  0.425000 2.495000 0.655000 ;
      RECT 2.325000  0.655000 3.505000 0.825000 ;
      RECT 2.325000  2.005000 2.575000 2.465000 ;
      RECT 2.765000  0.085000 3.095000 0.485000 ;
      RECT 3.335000  0.255000 3.505000 0.655000 ;
      RECT 3.335000  1.665000 3.505000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a311o_1
MACRO sky130_fd_sc_hd__a311o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.440000 0.605000 2.620000 0.995000 ;
        RECT 2.440000 0.995000 2.675000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895000 0.605000 2.165000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495000 0.995000 1.710000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895000 0.995000 3.235000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.695000 0.995000 4.005000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.295000 0.845000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.085000 0.345000 0.885000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 1.015000  0.085000 1.345000 0.465000 ;
      RECT 1.015000  0.655000 1.695000 0.825000 ;
      RECT 1.015000  0.825000 1.185000 1.495000 ;
      RECT 1.015000  1.495000 3.965000 1.665000 ;
      RECT 1.160000  1.835000 1.380000 2.635000 ;
      RECT 1.525000  0.255000 2.960000 0.425000 ;
      RECT 1.525000  0.425000 1.695000 0.655000 ;
      RECT 1.590000  1.835000 3.025000 2.005000 ;
      RECT 1.590000  2.005000 1.840000 2.465000 ;
      RECT 2.125000  2.255000 2.455000 2.635000 ;
      RECT 2.715000  2.005000 3.025000 2.465000 ;
      RECT 2.790000  0.425000 2.960000 0.655000 ;
      RECT 2.790000  0.655000 3.965000 0.825000 ;
      RECT 3.220000  0.085000 3.550000 0.485000 ;
      RECT 3.795000  0.255000 3.965000 0.655000 ;
      RECT 3.795000  1.665000 3.965000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__a311o_2
MACRO sky130_fd_sc_hd__a311o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.945000 1.075000 7.275000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.255000 1.075000 6.040000 1.285000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.515000 1.075000 4.945000 1.285000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 1.075000 1.505000 1.285000 ;
        RECT 1.060000 1.285000 1.255000 1.625000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 0.745000 0.350000 1.625000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.904000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195000 0.295000 2.545000 0.465000 ;
        RECT 2.295000 0.465000 2.465000 0.715000 ;
        RECT 2.295000 0.715000 3.305000 0.885000 ;
        RECT 2.715000 1.545000 3.885000 1.715000 ;
        RECT 2.910000 0.885000 3.105000 1.545000 ;
        RECT 3.055000 0.295000 3.385000 0.465000 ;
        RECT 3.135000 0.465000 3.305000 0.715000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.095000  0.085000 0.345000 0.565000 ;
      RECT 0.175000  1.795000 0.345000 2.295000 ;
      RECT 0.175000  2.295000 2.025000 2.465000 ;
      RECT 0.515000  0.295000 0.845000 0.465000 ;
      RECT 0.515000  1.955000 0.845000 2.125000 ;
      RECT 0.595000  0.465000 0.765000 0.715000 ;
      RECT 0.595000  0.715000 2.025000 0.885000 ;
      RECT 0.595000  0.885000 0.765000 1.955000 ;
      RECT 1.015000  0.085000 1.185000 0.545000 ;
      RECT 1.015000  1.795000 1.185000 2.295000 ;
      RECT 1.355000  0.295000 1.685000 0.465000 ;
      RECT 1.435000  0.465000 1.605000 0.715000 ;
      RECT 1.435000  1.455000 2.385000 1.625000 ;
      RECT 1.435000  1.625000 1.605000 2.125000 ;
      RECT 1.855000  0.085000 2.025000 0.545000 ;
      RECT 1.855000  0.885000 2.025000 1.075000 ;
      RECT 1.855000  1.075000 2.705000 1.245000 ;
      RECT 1.855000  1.795000 2.025000 2.295000 ;
      RECT 2.195000  1.625000 2.385000 1.915000 ;
      RECT 2.195000  1.915000 6.765000 2.085000 ;
      RECT 2.295000  2.255000 2.625000 2.635000 ;
      RECT 2.715000  0.085000 2.885000 0.545000 ;
      RECT 3.135000  2.255000 3.465000 2.635000 ;
      RECT 3.275000  1.075000 4.320000 1.245000 ;
      RECT 3.555000  0.085000 4.065000 0.545000 ;
      RECT 3.975000  2.255000 4.305000 2.635000 ;
      RECT 4.150000  1.245000 4.320000 1.455000 ;
      RECT 4.150000  1.455000 6.685000 1.625000 ;
      RECT 4.275000  0.295000 4.605000 0.465000 ;
      RECT 4.355000  0.465000 4.525000 0.715000 ;
      RECT 4.355000  0.715000 6.005000 0.885000 ;
      RECT 4.475000  1.795000 4.645000 1.915000 ;
      RECT 4.475000  2.085000 4.645000 2.465000 ;
      RECT 4.775000  0.085000 4.945000 0.545000 ;
      RECT 4.815000  2.255000 5.175000 2.635000 ;
      RECT 5.255000  0.255000 7.270000 0.425000 ;
      RECT 5.255000  0.425000 6.345000 0.465000 ;
      RECT 5.375000  1.795000 5.545000 1.915000 ;
      RECT 5.375000  2.085000 5.545000 2.465000 ;
      RECT 5.675000  0.645000 6.005000 0.715000 ;
      RECT 5.715000  2.255000 6.045000 2.635000 ;
      RECT 6.175000  0.465000 6.345000 0.885000 ;
      RECT 6.515000  0.645000 6.845000 0.825000 ;
      RECT 6.515000  0.825000 6.685000 1.455000 ;
      RECT 6.595000  1.795000 6.765000 1.915000 ;
      RECT 6.595000  2.085000 6.765000 2.465000 ;
      RECT 6.935000  0.425000 7.270000 0.500000 ;
      RECT 6.935000  1.795000 7.270000 2.635000 ;
      RECT 7.015000  0.500000 7.270000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__a311o_4
MACRO sky130_fd_sc_hd__a311oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 0.265000 1.365000 0.660000 ;
        RECT 1.195000 0.660000 1.365000 0.995000 ;
        RECT 1.195000 0.995000 1.455000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.600000 0.265000 0.795000 0.995000 ;
        RECT 0.600000 0.995000 1.025000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.420000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.710000 0.995000 1.935000 1.835000 ;
        RECT 1.710000 1.835000 2.230000 2.005000 ;
        RECT 1.950000 2.005000 2.230000 2.355000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 0.995000 2.685000 1.325000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.659750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 0.255000 1.705000 0.655000 ;
        RECT 1.535000 0.655000 2.650000 0.825000 ;
        RECT 2.105000 0.825000 2.275000 1.495000 ;
        RECT 2.105000 1.495000 2.650000 1.665000 ;
        RECT 2.405000 0.295000 2.650000 0.655000 ;
        RECT 2.410000 1.665000 2.650000 2.335000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.805000 ;
      RECT 0.095000  1.495000 0.425000 2.635000 ;
      RECT 0.600000  1.575000 1.540000 1.745000 ;
      RECT 0.600000  1.745000 0.770000 2.305000 ;
      RECT 0.940000  1.915000 1.200000 2.635000 ;
      RECT 1.370000  1.745000 1.540000 2.175000 ;
      RECT 1.370000  2.175000 1.700000 2.345000 ;
      RECT 1.905000  0.085000 2.235000 0.485000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a311oi_1
MACRO sky130_fd_sc_hd__a311oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.000000 0.995000 3.115000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 0.995000 1.805000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 0.995000 0.800000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395000 0.995000 4.055000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.730000 1.075000 5.410000 1.295000 ;
        RECT 5.175000 1.295000 5.410000 1.625000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.141000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295000 0.655000 5.345000 0.825000 ;
        RECT 3.235000 0.255000 3.405000 0.655000 ;
        RECT 4.085000 0.255000 4.255000 0.655000 ;
        RECT 4.260000 0.825000 4.475000 1.510000 ;
        RECT 4.260000 1.510000 4.990000 1.575000 ;
        RECT 4.260000 1.575000 5.005000 1.680000 ;
        RECT 4.660000 1.680000 5.005000 1.745000 ;
        RECT 4.660000 1.745000 4.990000 1.915000 ;
        RECT 4.660000 1.915000 5.005000 2.085000 ;
        RECT 5.175000 0.255000 5.345000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.095000  1.495000 0.345000 2.635000 ;
      RECT 0.175000  0.255000 0.345000 0.655000 ;
      RECT 0.175000  0.655000 2.105000 0.825000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.595000  1.575000 3.915000 1.745000 ;
      RECT 0.595000  1.745000 0.765000 2.465000 ;
      RECT 0.935000  1.915000 1.265000 2.635000 ;
      RECT 1.015000  0.255000 1.185000 0.655000 ;
      RECT 1.355000  0.305000 3.045000 0.475000 ;
      RECT 1.435000  1.745000 1.605000 2.465000 ;
      RECT 1.785000  1.915000 2.135000 2.635000 ;
      RECT 2.305000  1.745000 2.475000 2.465000 ;
      RECT 2.645000  1.915000 2.975000 2.635000 ;
      RECT 3.145000  2.255000 5.345000 2.425000 ;
      RECT 3.585000  0.085000 3.915000 0.465000 ;
      RECT 3.585000  1.745000 3.915000 2.085000 ;
      RECT 4.110000  1.915000 4.440000 2.255000 ;
      RECT 4.110000  2.425000 4.440000 2.465000 ;
      RECT 4.675000  0.085000 5.005000 0.465000 ;
      RECT 5.175000  1.795000 5.345000 2.255000 ;
      RECT 5.175000  2.425000 5.345000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__a311oi_2
MACRO sky130_fd_sc_hd__a311oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.995000 5.420000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.995000 3.550000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.995000 1.735000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.670000 0.995000 6.855000 1.630000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.935000 0.995000 9.530000 1.325000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.898500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.975000 0.635000 9.485000 0.805000 ;
        RECT 6.575000 0.255000 6.745000 0.635000 ;
        RECT 7.415000 0.255000 7.585000 0.635000 ;
        RECT 7.415000 0.805000 7.735000 1.545000 ;
        RECT 7.415000 1.545000 9.145000 1.715000 ;
        RECT 7.415000 1.715000 7.735000 1.975000 ;
        RECT 7.975000 1.530000 8.305000 1.545000 ;
        RECT 7.975000 1.715000 8.305000 2.085000 ;
        RECT 8.475000 0.255000 8.645000 0.635000 ;
        RECT 8.815000 1.715000 9.145000 2.085000 ;
        RECT 9.315000 0.255000 9.485000 0.635000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.095000  1.575000 0.425000 2.635000 ;
      RECT 0.175000  0.255000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 3.785000 0.805000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.595000  1.495000 4.965000 1.665000 ;
      RECT 0.595000  1.665000 0.765000 2.465000 ;
      RECT 0.935000  1.915000 1.265000 2.635000 ;
      RECT 1.015000  0.255000 1.185000 0.635000 ;
      RECT 1.355000  0.085000 1.685000 0.465000 ;
      RECT 1.435000  1.665000 1.605000 2.465000 ;
      RECT 1.775000  1.915000 2.105000 2.635000 ;
      RECT 1.855000  0.255000 2.025000 0.635000 ;
      RECT 2.195000  0.295000 5.565000 0.465000 ;
      RECT 2.275000  1.665000 2.445000 2.465000 ;
      RECT 2.615000  1.915000 2.945000 2.635000 ;
      RECT 3.115000  1.665000 3.285000 2.465000 ;
      RECT 3.455000  1.915000 3.785000 2.635000 ;
      RECT 3.955000  1.665000 4.125000 2.465000 ;
      RECT 4.295000  1.915000 4.625000 2.635000 ;
      RECT 4.795000  1.665000 4.965000 1.915000 ;
      RECT 4.795000  1.915000 7.245000 2.085000 ;
      RECT 4.795000  2.085000 4.965000 2.465000 ;
      RECT 5.135000  2.255000 5.465000 2.635000 ;
      RECT 5.655000  2.255000 9.565000 2.425000 ;
      RECT 6.075000  0.085000 6.405000 0.465000 ;
      RECT 6.915000  0.085000 7.245000 0.465000 ;
      RECT 7.975000  0.085000 8.305000 0.465000 ;
      RECT 8.815000  0.085000 9.145000 0.465000 ;
      RECT 9.315000  1.835000 9.565000 2.255000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
END sky130_fd_sc_hd__a311oi_4
MACRO sky130_fd_sc_hd__a2111o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.995000 3.290000 1.325000 ;
        RECT 2.985000 0.285000 3.540000 0.845000 ;
        RECT 2.985000 0.845000 3.290000 0.995000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.510000 1.025000 4.010000 1.290000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.400000 0.995000 2.680000 2.465000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.890000 1.050000 2.220000 2.465000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.290000 1.050000 1.720000 1.290000 ;
        RECT 1.515000 1.290000 1.720000 2.465000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.504500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 0.255000 0.465000 1.620000 ;
        RECT 0.135000 1.620000 0.390000 2.460000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
    PORT
      LAYER pwell ;
        RECT 1.975000 -0.065000 2.145000 0.105000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.565000  1.815000 0.895000 2.635000 ;
      RECT 0.635000  0.085000 1.310000 0.470000 ;
      RECT 0.695000  0.650000 1.915000 0.655000 ;
      RECT 0.695000  0.655000 2.805000 0.825000 ;
      RECT 0.695000  0.825000 0.915000 1.465000 ;
      RECT 0.695000  1.465000 1.345000 1.645000 ;
      RECT 1.135000  1.645000 1.345000 2.460000 ;
      RECT 1.585000  0.260000 1.915000 0.650000 ;
      RECT 2.085000  0.085000 2.430000 0.485000 ;
      RECT 2.600000  0.260000 2.805000 0.655000 ;
      RECT 2.860000  1.495000 3.990000 1.665000 ;
      RECT 2.860000  1.665000 3.145000 2.460000 ;
      RECT 3.325000  1.835000 3.540000 2.635000 ;
      RECT 3.715000  0.085000 3.955000 0.760000 ;
      RECT 3.720000  1.665000 3.990000 2.460000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__a2111o_1
MACRO sky130_fd_sc_hd__a2111o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 0.955000 3.775000 1.740000 ;
        RECT 3.505000 0.290000 3.995000 0.825000 ;
        RECT 3.505000 0.825000 3.775000 0.955000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.945000 0.995000 4.515000 1.740000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.995000 3.195000 1.740000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.425000 0.995000 2.735000 2.355000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885000 0.995000 2.255000 1.325000 ;
        RECT 1.960000 1.325000 2.255000 2.355000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.255000 0.895000 2.390000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.085000 0.435000 0.885000 ;
      RECT 0.085000  1.635000 0.435000 2.635000 ;
      RECT 1.065000  0.085000 2.010000 0.445000 ;
      RECT 1.065000  0.445000 1.325000 0.865000 ;
      RECT 1.065000  1.075000 1.705000 1.325000 ;
      RECT 1.065000  1.495000 1.315000 2.635000 ;
      RECT 1.495000  0.615000 3.335000 0.785000 ;
      RECT 1.495000  0.785000 1.705000 1.075000 ;
      RECT 1.495000  1.325000 1.705000 1.495000 ;
      RECT 1.495000  1.495000 1.785000 2.465000 ;
      RECT 2.180000  0.255000 2.420000 0.615000 ;
      RECT 2.590000  0.085000 2.920000 0.445000 ;
      RECT 3.070000  1.915000 4.515000 2.085000 ;
      RECT 3.070000  2.085000 3.400000 2.465000 ;
      RECT 3.090000  0.255000 3.335000 0.615000 ;
      RECT 3.590000  2.255000 3.920000 2.635000 ;
      RECT 4.090000  2.085000 4.515000 2.465000 ;
      RECT 4.165000  0.085000 4.515000 0.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__a2111o_2
MACRO sky130_fd_sc_hd__a2111o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825000 1.075000 4.495000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.675000 1.075000 5.625000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.450000 0.975000 3.255000 1.285000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.040000 0.975000 2.280000 1.285000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.370000 1.625000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.165000 0.255000 6.355000 0.635000 ;
        RECT 6.165000 0.635000 7.735000 0.805000 ;
        RECT 6.165000 1.465000 7.735000 1.635000 ;
        RECT 6.165000 1.635000 7.215000 1.715000 ;
        RECT 6.165000 1.715000 6.355000 2.465000 ;
        RECT 7.025000 0.255000 7.215000 0.635000 ;
        RECT 7.025000 1.715000 7.215000 2.465000 ;
        RECT 7.490000 0.805000 7.735000 1.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.110000  1.795000 0.370000 2.295000 ;
      RECT 0.110000  2.295000 2.160000 2.465000 ;
      RECT 0.180000  0.255000 0.440000 0.635000 ;
      RECT 0.180000  0.635000 3.655000 0.805000 ;
      RECT 0.540000  0.805000 0.870000 2.125000 ;
      RECT 0.610000  0.085000 0.940000 0.465000 ;
      RECT 1.040000  1.455000 1.230000 2.295000 ;
      RECT 1.110000  0.255000 1.340000 0.615000 ;
      RECT 1.110000  0.615000 3.655000 0.635000 ;
      RECT 1.400000  1.455000 3.100000 1.625000 ;
      RECT 1.400000  1.625000 1.730000 2.125000 ;
      RECT 1.510000  0.085000 1.840000 0.445000 ;
      RECT 1.900000  1.795000 2.160000 2.295000 ;
      RECT 2.015000  0.255000 2.240000 0.615000 ;
      RECT 2.340000  1.795000 2.675000 2.295000 ;
      RECT 2.340000  2.295000 3.650000 2.465000 ;
      RECT 2.420000  0.085000 3.295000 0.445000 ;
      RECT 2.845000  1.625000 3.100000 2.125000 ;
      RECT 3.320000  1.795000 5.495000 1.995000 ;
      RECT 3.320000  1.995000 3.650000 2.295000 ;
      RECT 3.465000  0.255000 4.585000 0.445000 ;
      RECT 3.465000  0.445000 3.655000 0.615000 ;
      RECT 3.465000  0.805000 3.655000 1.445000 ;
      RECT 3.465000  1.445000 5.975000 1.625000 ;
      RECT 3.825000  0.615000 5.495000 0.785000 ;
      RECT 3.865000  2.165000 4.195000 2.635000 ;
      RECT 4.365000  1.995000 4.625000 2.415000 ;
      RECT 4.805000  0.085000 5.140000 0.445000 ;
      RECT 4.805000  2.255000 5.140000 2.635000 ;
      RECT 5.310000  0.255000 5.495000 0.615000 ;
      RECT 5.310000  1.995000 5.495000 2.465000 ;
      RECT 5.665000  0.085000 5.995000 0.515000 ;
      RECT 5.665000  1.800000 5.995000 2.635000 ;
      RECT 5.795000  1.075000 7.320000 1.245000 ;
      RECT 5.795000  1.245000 5.975000 1.445000 ;
      RECT 6.525000  0.085000 6.855000 0.445000 ;
      RECT 6.525000  1.885000 6.855000 2.635000 ;
      RECT 7.385000  0.085000 7.715000 0.465000 ;
      RECT 7.385000  1.805000 7.715000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__a2111o_4
MACRO sky130_fd_sc_hd__a2111oi_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111oi_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.035000 1.070000 2.625000 1.400000 ;
        RECT 2.355000 0.660000 2.625000 1.070000 ;
        RECT 2.355000 1.400000 2.625000 1.735000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.795000 0.650000 3.135000 1.735000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495000 1.055000 1.845000 1.735000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 1.055000 1.325000 2.360000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.730000 0.435000 1.655000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  0.424000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.360000 1.825000 0.785000 2.465000 ;
        RECT 0.605000 0.635000 2.040000 0.885000 ;
        RECT 0.605000 0.885000 0.785000 1.825000 ;
        RECT 0.785000 0.255000 1.040000 0.615000 ;
        RECT 0.785000 0.615000 2.040000 0.635000 ;
        RECT 1.710000 0.280000 2.040000 0.615000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.285000  0.085000 0.615000 0.465000 ;
      RECT 1.210000  0.085000 1.540000 0.445000 ;
      RECT 1.540000  1.905000 2.870000 2.085000 ;
      RECT 1.540000  2.085000 1.870000 2.465000 ;
      RECT 2.040000  2.255000 2.370000 2.635000 ;
      RECT 2.470000  0.085000 2.800000 0.480000 ;
      RECT 2.540000  2.085000 2.870000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a2111oi_0
MACRO sky130_fd_sc_hd__a2111oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.440000 0.995000 2.725000 1.400000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.350000 3.090000 1.020000 ;
        RECT 2.905000 1.020000 3.540000 1.290000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.940000 1.050000 2.270000 1.400000 ;
        RECT 1.940000 1.400000 2.215000 2.455000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 1.050000 1.770000 2.455000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.785000 1.050000 1.235000 2.455000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.388750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.700000 1.375000 0.705000 ;
        RECT 0.145000 0.705000 2.420000 0.815000 ;
        RECT 0.145000 0.815000 2.300000 0.880000 ;
        RECT 0.145000 0.880000 0.530000 2.460000 ;
        RECT 1.045000 0.260000 1.375000 0.700000 ;
        RECT 2.090000 0.305000 2.420000 0.705000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
    PORT
      LAYER pwell ;
        RECT 1.975000 -0.065000 2.145000 0.105000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.315000  0.085000 0.630000 0.525000 ;
      RECT 1.550000  0.085000 1.880000 0.535000 ;
      RECT 2.395000  1.580000 3.505000 1.750000 ;
      RECT 2.395000  1.750000 2.625000 2.460000 ;
      RECT 2.800000  1.920000 3.130000 2.635000 ;
      RECT 3.270000  0.085000 3.510000 0.760000 ;
      RECT 3.310000  1.750000 3.505000 2.460000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a2111oi_1
MACRO sky130_fd_sc_hd__a2111oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.465000 0.985000 3.715000 1.445000 ;
        RECT 3.465000 1.445000 5.290000 1.675000 ;
        RECT 4.895000 0.995000 5.290000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.970000 1.015000 4.725000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.185000 1.030000 2.855000 1.275000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.045000 0.455000 1.445000 ;
        RECT 0.125000 1.445000 1.800000 1.680000 ;
        RECT 1.615000 1.030000 1.975000 1.275000 ;
        RECT 1.615000 1.275000 1.800000 1.445000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.755000 1.075000 1.425000 1.275000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.212750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.255000 0.380000 0.615000 ;
        RECT 0.120000 0.615000 5.355000 0.805000 ;
        RECT 0.120000 0.805000 3.255000 0.845000 ;
        RECT 0.900000 1.850000 2.140000 2.105000 ;
        RECT 1.050000 0.255000 1.295000 0.615000 ;
        RECT 1.965000 0.255000 2.295000 0.615000 ;
        RECT 1.970000 1.445000 3.255000 1.625000 ;
        RECT 1.970000 1.625000 2.140000 1.850000 ;
        RECT 2.965000 0.275000 3.295000 0.615000 ;
        RECT 3.025000 0.845000 3.255000 1.445000 ;
        RECT 5.020000 0.295000 5.355000 0.615000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.100000  1.870000 0.460000 2.275000 ;
      RECT 0.100000  2.275000 2.185000 2.295000 ;
      RECT 0.100000  2.295000 2.985000 2.465000 ;
      RECT 0.550000  0.085000 0.880000 0.445000 ;
      RECT 1.465000  0.085000 1.795000 0.445000 ;
      RECT 2.310000  1.795000 3.335000 1.845000 ;
      RECT 2.310000  1.845000 5.400000 1.965000 ;
      RECT 2.310000  1.965000 2.640000 2.060000 ;
      RECT 2.465000  0.085000 2.795000 0.445000 ;
      RECT 2.815000  2.135000 2.985000 2.295000 ;
      RECT 3.155000  1.965000 5.400000 2.095000 ;
      RECT 3.155000  2.095000 3.520000 2.465000 ;
      RECT 3.690000  2.275000 4.020000 2.635000 ;
      RECT 4.125000  0.085000 4.455000 0.445000 ;
      RECT 4.190000  2.095000 5.400000 2.105000 ;
      RECT 4.190000  2.105000 4.400000 2.465000 ;
      RECT 4.570000  2.275000 4.900000 2.635000 ;
      RECT 5.070000  2.105000 5.400000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__a2111oi_2
MACRO sky130_fd_sc_hd__a2111oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.095000 1.020000 7.745000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.960000 1.020000 9.990000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.955000 1.020000 5.650000 1.275000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.055000 1.020000 3.745000 1.275000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.495000 1.020000 1.845000 1.275000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  2.009500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.615000 7.620000 0.785000 ;
        RECT 0.145000 0.785000 0.320000 1.475000 ;
        RECT 0.145000 1.475000 1.720000 1.655000 ;
        RECT 0.530000 1.655000 1.720000 1.685000 ;
        RECT 0.530000 1.685000 0.860000 2.085000 ;
        RECT 0.615000 0.455000 0.790000 0.615000 ;
        RECT 1.390000 1.685000 1.720000 2.085000 ;
        RECT 1.460000 0.455000 1.650000 0.615000 ;
        RECT 2.400000 0.455000 2.590000 0.615000 ;
        RECT 3.260000 0.455000 3.510000 0.615000 ;
        RECT 4.180000 0.455000 4.420000 0.615000 ;
        RECT 5.090000 0.455000 5.275000 0.615000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.100000  1.835000  0.360000 2.255000 ;
      RECT 0.100000  2.255000  3.870000 2.445000 ;
      RECT 0.115000  0.085000  0.445000 0.445000 ;
      RECT 0.960000  0.085000  1.290000 0.445000 ;
      RECT 1.030000  1.855000  1.220000 2.255000 ;
      RECT 1.820000  0.085000  2.230000 0.445000 ;
      RECT 1.890000  1.855000  2.080000 2.255000 ;
      RECT 2.250000  1.475000  5.680000 1.655000 ;
      RECT 2.250000  1.655000  3.440000 1.685000 ;
      RECT 2.250000  1.685000  2.580000 2.085000 ;
      RECT 2.750000  1.855000  2.940000 2.255000 ;
      RECT 2.760000  0.085000  3.090000 0.445000 ;
      RECT 3.110000  1.685000  3.440000 2.085000 ;
      RECT 3.610000  1.835000  3.870000 2.255000 ;
      RECT 3.680000  0.085000  4.010000 0.445000 ;
      RECT 4.060000  1.835000  4.320000 2.255000 ;
      RECT 4.060000  2.255000  5.180000 2.275000 ;
      RECT 4.060000  2.275000  6.050000 2.445000 ;
      RECT 4.490000  1.655000  5.680000 1.685000 ;
      RECT 4.490000  1.685000  4.820000 2.085000 ;
      RECT 4.590000  0.085000  4.920000 0.445000 ;
      RECT 4.990000  1.855000  5.180000 2.255000 ;
      RECT 5.350000  1.685000  5.680000 2.085000 ;
      RECT 5.445000  0.085000  5.780000 0.445000 ;
      RECT 5.860000  1.445000  9.770000 1.615000 ;
      RECT 5.860000  1.615000  6.050000 2.275000 ;
      RECT 5.980000  0.275000  8.075000 0.445000 ;
      RECT 6.220000  1.785000  6.550000 2.635000 ;
      RECT 6.720000  1.615000  6.910000 2.315000 ;
      RECT 7.080000  1.805000  7.410000 2.635000 ;
      RECT 7.580000  1.615000  9.770000 1.665000 ;
      RECT 7.580000  1.665000  7.910000 2.315000 ;
      RECT 7.885000  0.445000  8.075000 0.615000 ;
      RECT 7.885000  0.615000  9.865000 0.785000 ;
      RECT 8.080000  1.895000  8.410000 2.635000 ;
      RECT 8.245000  0.085000  8.575000 0.445000 ;
      RECT 8.580000  1.665000  9.770000 1.670000 ;
      RECT 8.580000  1.670000  8.840000 2.290000 ;
      RECT 8.745000  0.300000  8.935000 0.615000 ;
      RECT 9.030000  1.915000  9.360000 2.635000 ;
      RECT 9.105000  0.085000  9.435000 0.445000 ;
      RECT 9.530000  1.670000  9.770000 2.260000 ;
      RECT 9.605000  0.290000  9.865000 0.615000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
END sky130_fd_sc_hd__a2111oi_4
MACRO sky130_fd_sc_hd__and2_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.185000 0.430000 1.955000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.940000 1.080000 1.270000 1.615000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.280900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.560000 0.255000 2.215000 0.525000 ;
        RECT 1.790000 1.835000 2.215000 2.465000 ;
        RECT 1.950000 0.525000 2.215000 1.835000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.160000  2.175000 0.430000 2.635000 ;
      RECT 0.185000  0.280000 0.490000 0.695000 ;
      RECT 0.185000  0.695000 1.780000 0.910000 ;
      RECT 0.185000  0.910000 0.770000 0.950000 ;
      RECT 0.600000  0.950000 0.770000 2.135000 ;
      RECT 0.600000  2.135000 0.865000 2.465000 ;
      RECT 0.950000  0.085000 1.390000 0.525000 ;
      RECT 1.110000  1.835000 1.620000 2.635000 ;
      RECT 1.450000  0.910000 1.780000 1.435000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__and2_0
MACRO sky130_fd_sc_hd__and2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.075000 0.775000 1.325000 ;
        RECT 0.100000 1.325000 0.365000 1.685000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 1.075000 1.335000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.657000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655000 0.255000 2.215000 0.545000 ;
        RECT 1.755000 1.915000 2.215000 2.465000 ;
        RECT 1.965000 0.545000 2.215000 1.915000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.285000  0.355000 0.615000 0.715000 ;
      RECT 0.285000  0.715000 1.675000 0.905000 ;
      RECT 0.285000  1.965000 0.565000 2.635000 ;
      RECT 0.735000  1.575000 1.675000 1.745000 ;
      RECT 0.735000  1.745000 1.035000 2.295000 ;
      RECT 1.235000  0.085000 1.485000 0.545000 ;
      RECT 1.235000  1.915000 1.565000 2.635000 ;
      RECT 1.505000  0.905000 1.675000 0.995000 ;
      RECT 1.505000  0.995000 1.795000 1.325000 ;
      RECT 1.505000  1.325000 1.675000 1.575000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__and2_1
MACRO sky130_fd_sc_hd__and2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.775000 1.325000 ;
        RECT 0.085000 1.325000 0.400000 1.765000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.075000 1.335000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.643500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.665000 0.255000 2.215000 0.545000 ;
        RECT 1.765000 1.915000 2.215000 2.465000 ;
        RECT 1.965000 0.545000 2.215000 1.915000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.285000  0.355000 0.615000 0.715000 ;
      RECT 0.285000  0.715000 1.675000 0.905000 ;
      RECT 0.285000  1.965000 0.565000 2.635000 ;
      RECT 0.735000  1.575000 1.675000 1.745000 ;
      RECT 0.735000  1.745000 1.035000 2.295000 ;
      RECT 1.245000  0.085000 1.495000 0.545000 ;
      RECT 1.245000  1.915000 1.575000 2.635000 ;
      RECT 1.505000  0.905000 1.675000 0.995000 ;
      RECT 1.505000  0.995000 1.795000 1.325000 ;
      RECT 1.505000  1.325000 1.675000 1.575000 ;
      RECT 2.385000  0.085000 2.675000 0.885000 ;
      RECT 2.385000  1.495000 2.675000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__and2_2
MACRO sky130_fd_sc_hd__and2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.995000 0.435000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.995000 0.980000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 0.515000 1.720000 0.615000 ;
        RECT 1.530000 0.615000 3.135000 0.845000 ;
        RECT 1.530000 1.535000 3.135000 1.760000 ;
        RECT 1.530000 1.760000 1.720000 2.465000 ;
        RECT 2.390000 0.255000 2.580000 0.615000 ;
        RECT 2.390000 1.760000 3.135000 1.765000 ;
        RECT 2.390000 1.765000 2.580000 2.465000 ;
        RECT 2.855000 0.845000 3.135000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.095000  0.255000 0.425000 0.615000 ;
      RECT 0.095000  0.615000 1.360000 0.805000 ;
      RECT 0.095000  1.880000 0.425000 2.635000 ;
      RECT 0.605000  1.580000 1.360000 1.750000 ;
      RECT 0.605000  1.750000 0.785000 2.465000 ;
      RECT 0.955000  0.085000 1.285000 0.445000 ;
      RECT 0.990000  1.935000 1.320000 2.635000 ;
      RECT 1.150000  0.805000 1.360000 1.020000 ;
      RECT 1.150000  1.020000 2.685000 1.355000 ;
      RECT 1.150000  1.355000 1.360000 1.580000 ;
      RECT 1.890000  0.085000 2.220000 0.445000 ;
      RECT 1.890000  1.935000 2.220000 2.635000 ;
      RECT 2.750000  0.085000 3.080000 0.445000 ;
      RECT 2.750000  1.935000 3.080000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__and2_4
MACRO sky130_fd_sc_hd__and2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.765000 0.445000 1.615000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 1.645000 2.175000 1.955000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.350000 1.580000 2.655000 2.365000 ;
        RECT 2.415000 0.255000 2.655000 0.775000 ;
        RECT 2.480000 0.775000 2.655000 1.580000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.590000 ;
      RECT 0.175000  1.785000 0.850000 2.015000 ;
      RECT 0.175000  2.015000 0.345000 2.445000 ;
      RECT 0.515000  2.185000 0.845000 2.635000 ;
      RECT 0.595000  0.280000 0.835000 0.655000 ;
      RECT 0.615000  0.655000 0.835000 0.805000 ;
      RECT 0.615000  0.805000 1.150000 1.135000 ;
      RECT 0.615000  1.135000 0.850000 1.785000 ;
      RECT 1.020000  1.305000 2.305000 1.325000 ;
      RECT 1.020000  1.325000 1.880000 1.475000 ;
      RECT 1.020000  1.475000 1.305000 2.420000 ;
      RECT 1.115000  0.270000 1.285000 0.415000 ;
      RECT 1.115000  0.415000 1.490000 0.610000 ;
      RECT 1.320000  0.610000 1.490000 0.945000 ;
      RECT 1.320000  0.945000 2.305000 1.305000 ;
      RECT 1.485000  2.165000 2.170000 2.635000 ;
      RECT 1.850000  0.085000 2.245000 0.580000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__and2b_1
MACRO sky130_fd_sc_hd__and2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.765000 0.450000 1.615000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.645000 2.200000 1.955000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 1.580000 2.680000 2.365000 ;
        RECT 2.445000 0.255000 2.680000 0.775000 ;
        RECT 2.505000 0.775000 2.680000 1.580000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.590000 ;
      RECT 0.175000  1.785000 0.855000 2.015000 ;
      RECT 0.175000  2.015000 0.345000 2.445000 ;
      RECT 0.515000  2.185000 0.845000 2.635000 ;
      RECT 0.595000  0.280000 0.835000 0.655000 ;
      RECT 0.620000  0.655000 0.835000 0.805000 ;
      RECT 0.620000  0.805000 1.175000 1.135000 ;
      RECT 0.620000  1.135000 0.855000 1.785000 ;
      RECT 1.045000  1.305000 2.335000 1.325000 ;
      RECT 1.045000  1.325000 1.905000 1.475000 ;
      RECT 1.045000  1.475000 1.330000 2.420000 ;
      RECT 1.115000  0.270000 1.285000 0.415000 ;
      RECT 1.115000  0.415000 1.515000 0.610000 ;
      RECT 1.345000  0.610000 1.515000 0.945000 ;
      RECT 1.345000  0.945000 2.335000 1.305000 ;
      RECT 1.510000  2.165000 2.195000 2.635000 ;
      RECT 1.875000  0.085000 2.275000 0.580000 ;
      RECT 2.865000  0.085000 3.135000 0.720000 ;
      RECT 2.865000  1.680000 3.135000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__and2b_2
MACRO sky130_fd_sc_hd__and2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.900000 0.625000 3.155000 0.995000 ;
        RECT 2.900000 0.995000 3.205000 1.325000 ;
        RECT 2.900000 1.325000 3.155000 1.745000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 0.995000 0.975000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.934000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.535000 2.730000 1.745000 ;
        RECT 1.525000 0.495000 1.715000 0.615000 ;
        RECT 1.525000 0.615000 2.730000 0.825000 ;
        RECT 2.440000 0.825000 2.730000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.615000 ;
      RECT 0.090000  0.615000 1.355000 0.805000 ;
      RECT 0.090000  2.255000 0.425000 2.635000 ;
      RECT 0.165000  0.995000 0.425000 1.325000 ;
      RECT 0.165000  1.325000 0.335000 1.915000 ;
      RECT 0.165000  1.915000 3.505000 2.085000 ;
      RECT 0.515000  1.500000 1.315000 1.745000 ;
      RECT 0.955000  0.085000 1.285000 0.445000 ;
      RECT 0.990000  2.275000 1.320000 2.635000 ;
      RECT 1.110000  1.435000 1.320000 1.485000 ;
      RECT 1.110000  1.485000 1.315000 1.500000 ;
      RECT 1.145000  0.805000 1.355000 0.995000 ;
      RECT 1.145000  0.995000 2.260000 1.355000 ;
      RECT 1.145000  1.355000 1.320000 1.435000 ;
      RECT 1.885000  0.085000 2.215000 0.445000 ;
      RECT 1.905000  2.275000 2.235000 2.635000 ;
      RECT 2.745000  0.085000 3.075000 0.445000 ;
      RECT 2.745000  2.275000 3.075000 2.635000 ;
      RECT 3.330000  0.495000 3.500000 0.675000 ;
      RECT 3.330000  0.675000 3.545000 0.845000 ;
      RECT 3.335000  1.530000 3.545000 1.700000 ;
      RECT 3.335000  1.700000 3.505000 1.915000 ;
      RECT 3.375000  0.845000 3.545000 1.530000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__and2b_4
MACRO sky130_fd_sc_hd__and3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.635000 0.635000 1.020000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 2.125000 1.345000 2.465000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.145000 0.305000 1.365000 0.790000 ;
        RECT 1.145000 0.790000 1.475000 1.215000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.940000 1.765000 2.215000 2.465000 ;
        RECT 1.955000 0.255000 2.215000 0.735000 ;
        RECT 2.045000 0.735000 2.215000 1.765000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.085000  0.295000 0.975000 0.465000 ;
      RECT 0.085000  1.190000 0.975000 1.260000 ;
      RECT 0.085000  1.260000 0.980000 1.285000 ;
      RECT 0.085000  1.285000 0.990000 1.300000 ;
      RECT 0.085000  1.300000 0.995000 1.315000 ;
      RECT 0.085000  1.315000 1.005000 1.320000 ;
      RECT 0.085000  1.320000 1.010000 1.330000 ;
      RECT 0.085000  1.330000 1.015000 1.340000 ;
      RECT 0.085000  1.340000 1.025000 1.345000 ;
      RECT 0.085000  1.345000 1.035000 1.355000 ;
      RECT 0.085000  1.355000 1.045000 1.360000 ;
      RECT 0.085000  1.360000 0.345000 1.810000 ;
      RECT 0.085000  1.980000 0.700000 2.080000 ;
      RECT 0.085000  2.080000 0.690000 2.635000 ;
      RECT 0.515000  1.710000 0.845000 1.955000 ;
      RECT 0.515000  1.955000 0.700000 1.980000 ;
      RECT 0.710000  1.360000 1.045000 1.365000 ;
      RECT 0.710000  1.365000 1.060000 1.370000 ;
      RECT 0.710000  1.370000 1.075000 1.380000 ;
      RECT 0.710000  1.380000 1.100000 1.385000 ;
      RECT 0.710000  1.385000 1.875000 1.390000 ;
      RECT 0.740000  1.390000 1.875000 1.425000 ;
      RECT 0.775000  1.425000 1.875000 1.450000 ;
      RECT 0.805000  0.465000 0.975000 1.190000 ;
      RECT 0.805000  1.450000 1.875000 1.480000 ;
      RECT 0.825000  1.480000 1.875000 1.510000 ;
      RECT 0.845000  1.510000 1.875000 1.540000 ;
      RECT 0.915000  1.540000 1.875000 1.550000 ;
      RECT 0.940000  1.550000 1.875000 1.560000 ;
      RECT 0.960000  1.560000 1.875000 1.575000 ;
      RECT 0.980000  1.575000 1.875000 1.590000 ;
      RECT 0.985000  1.590000 1.770000 1.600000 ;
      RECT 1.000000  1.600000 1.770000 1.635000 ;
      RECT 1.015000  1.635000 1.770000 1.885000 ;
      RECT 1.515000  2.090000 1.770000 2.635000 ;
      RECT 1.535000  0.085000 1.785000 0.625000 ;
      RECT 1.645000  0.990000 1.875000 1.385000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__and3_1
MACRO sky130_fd_sc_hd__and3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.470000 1.245000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.895000 2.125000 1.370000 2.465000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.305000 1.295000 0.750000 ;
        RECT 1.065000 0.750000 1.475000 1.245000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.970000 1.795000 2.245000 2.465000 ;
        RECT 1.980000 0.255000 2.230000 0.715000 ;
        RECT 2.060000 0.715000 2.230000 0.925000 ;
        RECT 2.060000 0.925000 2.675000 1.445000 ;
        RECT 2.075000 1.445000 2.245000 1.795000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  2.130000 0.715000 2.635000 ;
      RECT 0.100000  1.425000 1.890000 1.595000 ;
      RECT 0.100000  1.595000 0.355000 1.960000 ;
      RECT 0.105000  0.305000 0.895000 0.570000 ;
      RECT 0.525000  1.765000 0.855000 1.955000 ;
      RECT 0.525000  1.955000 0.715000 2.130000 ;
      RECT 0.640000  0.570000 0.895000 1.425000 ;
      RECT 1.080000  1.595000 1.330000 1.890000 ;
      RECT 1.475000  0.085000 1.805000 0.580000 ;
      RECT 1.555000  1.790000 1.770000 2.635000 ;
      RECT 1.660000  0.995000 1.890000 1.425000 ;
      RECT 2.400000  0.085000 2.675000 0.745000 ;
      RECT 2.415000  1.625000 2.675000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__and3_2
MACRO sky130_fd_sc_hd__and3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.995000 0.875000 1.340000 ;
        RECT 0.115000 1.340000 0.365000 2.335000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.745000 1.355000 1.340000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.995000 1.900000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.450000 0.515000 2.640000 0.615000 ;
        RECT 2.450000 0.615000 4.055000 0.845000 ;
        RECT 2.450000 1.535000 4.055000 1.760000 ;
        RECT 2.450000 1.760000 2.640000 2.465000 ;
        RECT 3.310000 0.255000 3.500000 0.615000 ;
        RECT 3.310000 1.760000 4.055000 1.765000 ;
        RECT 3.310000 1.765000 3.500000 2.465000 ;
        RECT 3.775000 0.845000 4.055000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.465000  0.255000 0.800000 0.375000 ;
      RECT 0.465000  0.375000 1.725000 0.565000 ;
      RECT 0.465000  0.565000 0.800000 0.805000 ;
      RECT 0.545000  1.580000 2.280000 1.750000 ;
      RECT 0.545000  1.750000 0.725000 2.465000 ;
      RECT 0.895000  1.935000 1.345000 2.635000 ;
      RECT 1.520000  1.750000 1.700000 2.465000 ;
      RECT 1.535000  0.565000 1.725000 0.615000 ;
      RECT 1.535000  0.615000 2.280000 0.805000 ;
      RECT 1.905000  0.085000 2.235000 0.445000 ;
      RECT 1.910000  1.935000 2.240000 2.635000 ;
      RECT 2.070000  0.805000 2.280000 1.020000 ;
      RECT 2.070000  1.020000 3.605000 1.355000 ;
      RECT 2.070000  1.355000 2.280000 1.580000 ;
      RECT 2.810000  0.085000 3.140000 0.445000 ;
      RECT 2.810000  1.935000 3.140000 2.635000 ;
      RECT 3.670000  0.085000 4.000000 0.445000 ;
      RECT 3.670000  1.935000 4.000000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__and3_4
MACRO sky130_fd_sc_hd__and3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.955000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.790000 2.125000 2.265000 2.465000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.305000 2.185000 0.725000 ;
        RECT 1.985000 0.725000 2.395000 1.245000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.860000 1.765000 3.135000 2.465000 ;
        RECT 2.875000 0.255000 3.135000 0.735000 ;
        RECT 2.965000 0.735000 3.135000 1.765000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.905000 ;
      RECT 0.085000  2.125000 0.345000 2.635000 ;
      RECT 0.515000  0.485000 0.845000 0.905000 ;
      RECT 0.595000  0.905000 0.845000 0.995000 ;
      RECT 0.595000  0.995000 1.390000 1.245000 ;
      RECT 0.595000  1.245000 0.765000 2.465000 ;
      RECT 1.005000  1.425000 2.795000 1.595000 ;
      RECT 1.005000  1.595000 1.255000 1.960000 ;
      RECT 1.005000  2.130000 1.620000 2.635000 ;
      RECT 1.025000  0.305000 1.815000 0.570000 ;
      RECT 1.425000  1.765000 1.755000 1.955000 ;
      RECT 1.425000  1.955000 1.620000 2.130000 ;
      RECT 1.560000  0.570000 1.815000 1.425000 ;
      RECT 1.975000  1.595000 2.690000 1.890000 ;
      RECT 2.375000  0.085000 2.705000 0.545000 ;
      RECT 2.435000  2.090000 2.650000 2.635000 ;
      RECT 2.565000  0.995000 2.795000 1.425000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__and3b_1
MACRO sky130_fd_sc_hd__and3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.745000 0.410000 1.325000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.815000 2.125000 2.290000 2.465000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.010000 0.305000 2.220000 0.765000 ;
        RECT 2.010000 0.765000 2.420000 1.245000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875000 1.795000 3.160000 2.465000 ;
        RECT 2.915000 0.255000 3.160000 0.715000 ;
        RECT 2.990000 0.715000 3.160000 0.925000 ;
        RECT 2.990000 0.925000 3.595000 1.445000 ;
        RECT 2.990000 1.445000 3.160000 1.795000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.085000 0.355000 0.575000 ;
      RECT 0.085000  1.575000 0.400000 2.635000 ;
      RECT 0.580000  0.305000 0.855000 1.015000 ;
      RECT 0.580000  1.015000 1.415000 1.245000 ;
      RECT 0.580000  1.245000 0.855000 1.905000 ;
      RECT 1.030000  2.130000 1.645000 2.635000 ;
      RECT 1.050000  1.425000 2.820000 1.595000 ;
      RECT 1.050000  1.595000 1.285000 1.960000 ;
      RECT 1.055000  0.305000 1.840000 0.570000 ;
      RECT 1.455000  1.765000 1.785000 1.955000 ;
      RECT 1.455000  1.955000 1.645000 2.130000 ;
      RECT 1.585000  0.570000 1.840000 1.425000 ;
      RECT 2.010000  1.595000 2.200000 1.890000 ;
      RECT 2.410000  0.085000 2.740000 0.580000 ;
      RECT 2.460000  1.790000 2.675000 2.635000 ;
      RECT 2.590000  0.995000 2.820000 1.425000 ;
      RECT 3.330000  0.085000 3.595000 0.745000 ;
      RECT 3.330000  1.625000 3.595000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__and3b_2
MACRO sky130_fd_sc_hd__and3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.715000 0.615000 3.995000 1.705000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.020000 0.725000 1.235000 1.340000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.995000 1.715000 1.340000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.934000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.225000 1.535000 3.535000 1.705000 ;
        RECT 2.285000 0.515000 2.475000 0.615000 ;
        RECT 2.285000 0.615000 3.535000 0.845000 ;
        RECT 3.145000 0.255000 3.335000 0.615000 ;
        RECT 3.270000 0.845000 3.535000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.150000  0.255000 0.635000 0.355000 ;
      RECT 0.150000  0.355000 1.600000 0.545000 ;
      RECT 0.150000  0.545000 0.635000 0.805000 ;
      RECT 0.150000  0.805000 0.370000 1.495000 ;
      RECT 0.150000  1.495000 0.510000 2.165000 ;
      RECT 0.540000  0.995000 0.850000 1.325000 ;
      RECT 0.680000  1.325000 0.850000 1.875000 ;
      RECT 0.680000  1.875000 4.445000 2.105000 ;
      RECT 0.730000  2.275000 1.180000 2.635000 ;
      RECT 1.280000  1.525000 2.055000 1.695000 ;
      RECT 1.420000  0.545000 1.600000 0.615000 ;
      RECT 1.420000  0.615000 2.115000 0.805000 ;
      RECT 1.745000  2.275000 2.075000 2.635000 ;
      RECT 1.780000  0.085000 2.110000 0.445000 ;
      RECT 1.885000  0.805000 2.115000 1.020000 ;
      RECT 1.885000  1.020000 3.100000 1.355000 ;
      RECT 1.885000  1.355000 2.055000 1.525000 ;
      RECT 2.645000  0.085000 2.975000 0.445000 ;
      RECT 2.645000  2.275000 2.980000 2.635000 ;
      RECT 3.505000  0.085000 3.835000 0.445000 ;
      RECT 3.505000  2.275000 3.835000 2.635000 ;
      RECT 4.165000  0.425000 4.445000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__and3b_4
MACRO sky130_fd_sc_hd__and4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.325000 2.075000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.885000 0.360000 1.235000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 0.355000 1.715000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895000 0.355000 2.175000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.795000 0.295000 3.135000 0.805000 ;
        RECT 2.795000 2.205000 3.135000 2.465000 ;
        RECT 2.875000 0.805000 3.135000 2.205000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  2.255000 0.425000 2.635000 ;
      RECT 0.170000  0.255000 0.665000 0.585000 ;
      RECT 0.495000  0.585000 0.665000 1.495000 ;
      RECT 0.495000  1.495000 2.685000 1.665000 ;
      RECT 0.595000  1.665000 0.845000 2.465000 ;
      RECT 1.065000  1.915000 1.395000 2.635000 ;
      RECT 1.580000  1.665000 1.830000 2.465000 ;
      RECT 2.295000  1.835000 2.625000 2.635000 ;
      RECT 2.355000  0.085000 2.625000 0.885000 ;
      RECT 2.370000  1.075000 2.700000 1.325000 ;
      RECT 2.370000  1.325000 2.685000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__and4_1
MACRO sky130_fd_sc_hd__and4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.755000 0.330000 2.075000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.890000 0.420000 1.245000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.420000 0.415000 1.720000 1.305000 ;
        RECT 1.420000 1.305000 1.590000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.900000 0.415000 2.160000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.544500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 0.295000 3.065000 0.340000 ;
        RECT 2.735000 0.340000 3.070000 0.805000 ;
        RECT 2.735000 1.495000 3.070000 2.465000 ;
        RECT 2.895000 0.805000 3.070000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.095000  2.255000 0.425000 2.635000 ;
      RECT 0.175000  0.255000 0.670000 0.585000 ;
      RECT 0.500000  0.585000 0.670000 1.495000 ;
      RECT 0.500000  1.495000 2.555000 1.665000 ;
      RECT 0.600000  1.665000 0.850000 2.465000 ;
      RECT 1.070000  1.915000 1.400000 2.635000 ;
      RECT 1.585000  1.665000 1.835000 2.465000 ;
      RECT 2.235000  1.835000 2.565000 2.635000 ;
      RECT 2.330000  0.085000 2.565000 0.890000 ;
      RECT 2.330000  1.075000 2.725000 1.315000 ;
      RECT 2.330000  1.315000 2.555000 1.495000 ;
      RECT 3.245000  1.835000 3.575000 2.635000 ;
      RECT 3.255000  0.085000 3.585000 0.810000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__and4_2
MACRO sky130_fd_sc_hd__and4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.765000 0.330000 1.655000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.840000 0.995000 1.245000 1.325000 ;
        RECT 0.890000 0.420000 1.245000 0.995000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 0.425000 1.700000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.905000 0.730000 2.155000 0.935000 ;
        RECT 1.905000 0.935000 2.075000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.535000 0.255000 2.705000 0.640000 ;
        RECT 2.535000 0.640000 4.050000 0.810000 ;
        RECT 2.535000 1.795000 2.785000 2.465000 ;
        RECT 2.615000 1.485000 4.050000 1.655000 ;
        RECT 2.615000 1.655000 2.785000 1.795000 ;
        RECT 3.375000 0.255000 3.545000 0.640000 ;
        RECT 3.375000 1.655000 4.050000 1.745000 ;
        RECT 3.375000 1.745000 3.545000 2.465000 ;
        RECT 3.800000 0.810000 4.050000 1.485000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.105000  1.835000 0.385000 2.635000 ;
      RECT 0.175000  0.255000 0.670000 0.585000 ;
      RECT 0.500000  0.585000 0.670000 1.495000 ;
      RECT 0.500000  1.495000 2.415000 1.665000 ;
      RECT 0.555000  1.665000 0.765000 2.465000 ;
      RECT 0.955000  1.935000 1.285000 2.635000 ;
      RECT 1.455000  1.665000 1.645000 2.465000 ;
      RECT 2.025000  0.085000 2.335000 0.550000 ;
      RECT 2.025000  1.855000 2.355000 2.635000 ;
      RECT 2.245000  1.105000 3.585000 1.305000 ;
      RECT 2.245000  1.305000 2.415000 1.495000 ;
      RECT 2.575000  1.075000 3.585000 1.105000 ;
      RECT 2.875000  0.085000 3.205000 0.470000 ;
      RECT 2.955000  1.835000 3.205000 2.635000 ;
      RECT 3.715000  0.085000 4.045000 0.470000 ;
      RECT 3.715000  1.915000 4.045000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__and4_4
MACRO sky130_fd_sc_hd__and4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.450000 1.675000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.520000 0.420000 1.800000 1.695000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025000 0.420000 2.295000 1.695000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485000 0.665000 2.825000 1.695000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.255000 0.295000 3.590000 0.340000 ;
        RECT 3.255000 0.340000 3.595000 0.805000 ;
        RECT 3.335000 1.495000 3.595000 2.465000 ;
        RECT 3.425000 0.805000 3.595000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.170000  0.255000 0.345000 0.655000 ;
      RECT 0.170000  0.655000 0.800000 0.825000 ;
      RECT 0.170000  1.845000 0.800000 2.015000 ;
      RECT 0.170000  2.015000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.195000 0.845000 2.635000 ;
      RECT 0.630000  0.825000 0.800000 0.995000 ;
      RECT 0.630000  0.995000 0.980000 1.325000 ;
      RECT 0.630000  1.325000 0.800000 1.845000 ;
      RECT 1.090000  0.255000 1.320000 0.585000 ;
      RECT 1.150000  0.585000 1.320000 1.875000 ;
      RECT 1.150000  1.875000 3.165000 2.045000 ;
      RECT 1.150000  2.045000 1.320000 2.465000 ;
      RECT 1.555000  2.225000 2.225000 2.635000 ;
      RECT 2.440000  2.045000 2.610000 2.465000 ;
      RECT 2.755000  0.085000 3.085000 0.465000 ;
      RECT 2.810000  2.225000 3.140000 2.635000 ;
      RECT 2.995000  0.995000 3.255000 1.325000 ;
      RECT 2.995000  1.325000 3.165000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__and4b_1
MACRO sky130_fd_sc_hd__and4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 0.740000 0.335000 1.630000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.420000 1.745000 1.745000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.960000 0.420000 2.275000 1.695000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 0.645000 2.775000 1.615000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.503250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.260000 0.255000 3.545000 0.640000 ;
        RECT 3.260000 0.640000 4.055000 0.825000 ;
        RECT 3.340000 1.535000 4.055000 1.745000 ;
        RECT 3.340000 1.745000 3.545000 2.465000 ;
        RECT 3.425000 0.825000 4.055000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.175000  1.830000 0.805000 2.000000 ;
      RECT 0.175000  2.000000 0.345000 2.465000 ;
      RECT 0.515000  2.195000 0.845000 2.635000 ;
      RECT 0.595000  0.255000 0.805000 0.585000 ;
      RECT 0.635000  0.585000 0.805000 0.995000 ;
      RECT 0.635000  0.995000 0.975000 1.325000 ;
      RECT 0.635000  1.325000 0.805000 1.830000 ;
      RECT 1.015000  1.660000 1.315000 1.915000 ;
      RECT 1.015000  1.915000 3.165000 1.965000 ;
      RECT 1.015000  1.965000 2.610000 2.085000 ;
      RECT 1.015000  2.085000 1.185000 2.465000 ;
      RECT 1.095000  0.255000 1.315000 0.585000 ;
      RECT 1.145000  0.585000 1.315000 1.660000 ;
      RECT 1.555000  2.255000 2.225000 2.635000 ;
      RECT 2.440000  1.795000 3.165000 1.915000 ;
      RECT 2.440000  2.085000 2.610000 2.465000 ;
      RECT 2.760000  0.085000 3.090000 0.465000 ;
      RECT 2.840000  2.195000 3.170000 2.635000 ;
      RECT 2.995000  0.995000 3.255000 1.325000 ;
      RECT 2.995000  1.325000 3.165000 1.795000 ;
      RECT 3.715000  0.085000 4.050000 0.465000 ;
      RECT 3.715000  1.915000 4.050000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__and4b_2
MACRO sky130_fd_sc_hd__and4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 0.765000 0.790000 1.635000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 0.735000 4.145000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.345000 0.755000 3.555000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865000 0.995000 3.085000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.980000 0.650000 2.080000 0.820000 ;
        RECT 0.980000 0.820000 1.260000 1.545000 ;
        RECT 0.980000 1.545000 2.160000 1.715000 ;
        RECT 1.070000 0.255000 1.240000 0.650000 ;
        RECT 1.910000 0.255000 2.080000 0.650000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.585000 ;
      RECT 0.085000  0.585000 0.260000 1.915000 ;
      RECT 0.085000  1.915000 4.900000 2.085000 ;
      RECT 0.085000  2.085000 0.345000 2.465000 ;
      RECT 0.515000  2.255000 0.845000 2.635000 ;
      RECT 0.570000  0.085000 0.900000 0.470000 ;
      RECT 1.410000  0.085000 1.740000 0.470000 ;
      RECT 1.410000  2.255000 1.740000 2.635000 ;
      RECT 1.440000  1.075000 2.550000 1.245000 ;
      RECT 2.250000  2.255000 2.580000 2.635000 ;
      RECT 2.285000  0.085000 2.615000 0.445000 ;
      RECT 2.380000  0.615000 2.965000 0.785000 ;
      RECT 2.380000  0.785000 2.550000 1.075000 ;
      RECT 2.380000  1.245000 2.550000 1.545000 ;
      RECT 2.380000  1.545000 4.545000 1.715000 ;
      RECT 2.795000  0.300000 4.965000 0.470000 ;
      RECT 2.795000  0.470000 2.965000 0.615000 ;
      RECT 3.475000  2.255000 3.805000 2.635000 ;
      RECT 4.390000  0.470000 4.965000 0.810000 ;
      RECT 4.635000  2.255000 4.965000 2.635000 ;
      RECT 4.730000  0.995000 4.900000 1.915000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__and4b_4
MACRO sky130_fd_sc_hd__and4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.625000 0.775000 1.955000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.765000 0.815000 0.945000 ;
        RECT 0.605000 0.945000 1.225000 1.115000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895000 0.415000 3.080000 0.995000 ;
        RECT 2.895000 0.995000 3.125000 1.325000 ;
        RECT 2.895000 1.325000 3.080000 1.635000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.350000 0.420000 3.545000 0.995000 ;
        RECT 3.350000 0.995000 3.605000 1.325000 ;
        RECT 3.350000 1.325000 3.545000 1.635000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.425400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.255000 0.255000 4.515000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.585000 ;
      RECT 0.085000  0.585000 0.255000 1.285000 ;
      RECT 0.085000  1.285000 1.215000 1.455000 ;
      RECT 0.085000  1.455000 0.255000 2.135000 ;
      RECT 0.085000  2.135000 0.345000 2.465000 ;
      RECT 0.655000  0.085000 0.985000 0.465000 ;
      RECT 0.655000  2.255000 0.985000 2.635000 ;
      RECT 1.045000  1.455000 1.215000 1.575000 ;
      RECT 1.045000  1.575000 1.625000 1.745000 ;
      RECT 1.165000  0.255000 2.645000 0.425000 ;
      RECT 1.165000  0.425000 1.565000 0.755000 ;
      RECT 1.225000  1.915000 1.965000 2.085000 ;
      RECT 1.225000  2.085000 1.415000 2.465000 ;
      RECT 1.395000  0.755000 1.565000 1.235000 ;
      RECT 1.395000  1.235000 1.965000 1.405000 ;
      RECT 1.665000  2.255000 1.995000 2.635000 ;
      RECT 1.755000  0.595000 2.305000 0.925000 ;
      RECT 1.795000  1.405000 1.965000 1.915000 ;
      RECT 2.135000  0.925000 2.305000 1.915000 ;
      RECT 2.135000  1.915000 4.085000 2.085000 ;
      RECT 2.205000  2.085000 2.375000 2.465000 ;
      RECT 2.475000  0.425000 2.645000 1.325000 ;
      RECT 2.570000  2.255000 2.900000 2.635000 ;
      RECT 3.160000  2.085000 3.330000 2.465000 ;
      RECT 3.755000  0.085000 4.085000 0.465000 ;
      RECT 3.755000  2.255000 4.085000 2.635000 ;
      RECT 3.915000  0.995000 4.085000 1.915000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__and4bb_1
MACRO sky130_fd_sc_hd__and4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.995000 0.330000 1.635000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825000 0.765000 4.175000 1.305000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.910000 0.420000 3.175000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.350000 0.425000 3.655000 1.405000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.990000 1.545000 1.320000 1.715000 ;
        RECT 1.015000 0.255000 1.240000 1.545000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.175000  0.255000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.670000 0.805000 ;
      RECT 0.175000  1.885000 1.925000 2.055000 ;
      RECT 0.175000  2.055000 0.345000 2.465000 ;
      RECT 0.500000  0.805000 0.670000 1.885000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.255000 0.845000 2.635000 ;
      RECT 1.410000  0.085000 1.740000 0.465000 ;
      RECT 1.415000  0.635000 2.405000 0.805000 ;
      RECT 1.415000  0.805000 1.585000 1.325000 ;
      RECT 1.490000  2.255000 2.160000 2.635000 ;
      RECT 1.755000  0.995000 2.065000 1.325000 ;
      RECT 1.755000  1.325000 1.925000 1.885000 ;
      RECT 2.010000  0.255000 2.180000 0.635000 ;
      RECT 2.235000  0.805000 2.405000 1.915000 ;
      RECT 2.235000  1.915000 3.415000 2.085000 ;
      RECT 2.395000  2.085000 2.565000 2.465000 ;
      RECT 2.575000  1.400000 2.745000 1.575000 ;
      RECT 2.575000  1.575000 3.755000 1.745000 ;
      RECT 2.735000  2.255000 3.075000 2.635000 ;
      RECT 3.245000  2.085000 3.415000 2.465000 ;
      RECT 3.585000  1.745000 3.755000 1.915000 ;
      RECT 3.585000  1.915000 4.515000 2.085000 ;
      RECT 3.755000  2.255000 4.085000 2.635000 ;
      RECT 3.835000  0.085000 4.085000 0.585000 ;
      RECT 4.255000  0.255000 4.515000 0.585000 ;
      RECT 4.255000  2.085000 4.515000 2.465000 ;
      RECT 4.345000  0.585000 4.515000 1.915000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__and4bb_2
MACRO sky130_fd_sc_hd__and4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.485000 0.995000 5.845000 1.620000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.765000 0.780000 1.635000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.250000 0.755000 3.545000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.680000 0.995000 3.080000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.960000 0.650000 2.080000 0.820000 ;
        RECT 0.960000 0.820000 1.240000 1.545000 ;
        RECT 0.960000 1.545000 2.160000 1.715000 ;
        RECT 1.070000 0.255000 1.240000 0.650000 ;
        RECT 1.910000 0.255000 2.080000 0.650000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.585000 ;
      RECT 0.085000  0.585000 0.260000 1.915000 ;
      RECT 0.085000  1.915000 4.490000 2.085000 ;
      RECT 0.085000  2.085000 0.345000 2.465000 ;
      RECT 0.515000  2.255000 0.845000 2.635000 ;
      RECT 0.570000  0.085000 0.900000 0.470000 ;
      RECT 1.410000  0.085000 1.740000 0.470000 ;
      RECT 1.410000  1.075000 2.500000 1.245000 ;
      RECT 1.410000  2.255000 1.740000 2.635000 ;
      RECT 2.250000  2.255000 2.580000 2.635000 ;
      RECT 2.270000  0.085000 2.600000 0.445000 ;
      RECT 2.330000  0.615000 2.940000 0.785000 ;
      RECT 2.330000  0.785000 2.500000 1.075000 ;
      RECT 2.330000  1.245000 2.500000 1.545000 ;
      RECT 2.330000  1.545000 4.150000 1.715000 ;
      RECT 2.770000  0.300000 4.610000 0.470000 ;
      RECT 2.770000  0.470000 2.940000 0.615000 ;
      RECT 3.330000  2.255000 3.660000 2.635000 ;
      RECT 3.730000  0.995000 3.900000 1.155000 ;
      RECT 3.730000  1.155000 4.490000 1.325000 ;
      RECT 4.255000  0.470000 4.610000 0.810000 ;
      RECT 4.320000  1.325000 4.490000 1.915000 ;
      RECT 4.360000  2.255000 5.370000 2.635000 ;
      RECT 4.950000  0.655000 5.805000 0.825000 ;
      RECT 4.950000  0.825000 5.120000 1.915000 ;
      RECT 4.950000  1.915000 5.805000 2.085000 ;
      RECT 4.975000  0.085000 5.305000 0.465000 ;
      RECT 5.635000  0.255000 5.805000 0.655000 ;
      RECT 5.635000  2.085000 5.805000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__and4bb_4
MACRO sky130_fd_sc_hd__buf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.196500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.985000 0.445000 1.355000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 1.560000 1.295000 2.465000 ;
        RECT 1.035000 0.255000 1.295000 0.760000 ;
        RECT 1.115000 0.760000 1.295000 1.560000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.165000  1.535000 0.840000 1.705000 ;
      RECT 0.165000  1.705000 0.345000 2.465000 ;
      RECT 0.175000  0.255000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.840000 0.805000 ;
      RECT 0.525000  0.085000 0.855000 0.465000 ;
      RECT 0.525000  1.875000 0.855000 2.635000 ;
      RECT 0.670000  0.805000 0.840000 1.060000 ;
      RECT 0.670000  1.060000 0.945000 1.390000 ;
      RECT 0.670000  1.390000 0.840000 1.535000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__buf_1
MACRO sky130_fd_sc_hd__buf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.440000 1.355000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 0.255000 1.315000 0.830000 ;
        RECT 1.060000 1.560000 1.315000 2.465000 ;
        RECT 1.145000 0.830000 1.315000 1.560000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.175000  0.255000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.890000 0.805000 ;
      RECT 0.175000  1.535000 0.890000 1.705000 ;
      RECT 0.175000  1.705000 0.345000 2.465000 ;
      RECT 0.560000  0.085000 0.890000 0.465000 ;
      RECT 0.560000  1.875000 0.890000 2.635000 ;
      RECT 0.720000  0.805000 0.890000 0.995000 ;
      RECT 0.720000  0.995000 0.975000 1.325000 ;
      RECT 0.720000  1.325000 0.890000 1.535000 ;
      RECT 1.490000  0.085000 1.750000 0.925000 ;
      RECT 1.490000  1.485000 1.750000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__buf_2
MACRO sky130_fd_sc_hd__buf_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.470000 1.315000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 0.255000 1.185000 0.735000 ;
        RECT 1.015000 0.735000 2.025000 0.905000 ;
        RECT 1.015000 1.445000 2.025000 1.615000 ;
        RECT 1.015000 1.615000 1.185000 2.465000 ;
        RECT 1.530000 0.905000 2.025000 1.445000 ;
        RECT 1.855000 0.255000 2.025000 0.735000 ;
        RECT 1.855000 1.615000 2.025000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.095000  1.485000 0.810000 1.655000 ;
      RECT 0.095000  1.655000 0.425000 2.465000 ;
      RECT 0.175000  0.255000 0.345000 0.735000 ;
      RECT 0.175000  0.735000 0.810000 0.905000 ;
      RECT 0.525000  0.085000 0.765000 0.565000 ;
      RECT 0.595000  1.835000 0.835000 2.635000 ;
      RECT 0.640000  0.905000 0.810000 1.075000 ;
      RECT 0.640000  1.075000 1.140000 1.245000 ;
      RECT 0.640000  1.245000 0.810000 1.485000 ;
      RECT 1.355000  0.085000 1.685000 0.565000 ;
      RECT 1.355000  1.835000 1.685000 2.635000 ;
      RECT 2.195000  0.085000 2.525000 0.885000 ;
      RECT 2.195000  1.485000 2.525000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__buf_4
MACRO sky130_fd_sc_hd__buf_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_6 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.280000 1.075000 1.185000 1.315000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.336500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.255000 1.865000 0.735000 ;
        RECT 1.695000 0.735000 3.545000 0.905000 ;
        RECT 1.695000 1.445000 3.545000 1.615000 ;
        RECT 1.695000 1.615000 1.865000 2.465000 ;
        RECT 2.210000 0.905000 3.545000 1.445000 ;
        RECT 2.535000 0.255000 2.705000 0.735000 ;
        RECT 2.535000 1.615000 2.705000 2.465000 ;
        RECT 3.375000 0.255000 3.545000 0.735000 ;
        RECT 3.375000 1.615000 3.545000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.435000  0.085000 0.605000 0.565000 ;
      RECT 0.435000  1.485000 0.605000 2.635000 ;
      RECT 0.775000  0.255000 1.105000 0.735000 ;
      RECT 0.775000  0.735000 1.525000 0.905000 ;
      RECT 0.775000  1.485000 1.525000 1.655000 ;
      RECT 0.775000  1.655000 1.105000 2.465000 ;
      RECT 1.275000  0.085000 1.445000 0.565000 ;
      RECT 1.275000  1.835000 1.515000 2.635000 ;
      RECT 1.355000  0.905000 1.525000 1.075000 ;
      RECT 1.355000  1.075000 1.825000 1.245000 ;
      RECT 1.355000  1.245000 1.525000 1.485000 ;
      RECT 2.035000  0.085000 2.365000 0.565000 ;
      RECT 2.035000  1.835000 2.365000 2.635000 ;
      RECT 2.875000  0.085000 3.205000 0.565000 ;
      RECT 2.875000  1.835000 3.205000 2.635000 ;
      RECT 3.715000  0.085000 4.045000 0.885000 ;
      RECT 3.715000  1.485000 4.045000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__buf_6
MACRO sky130_fd_sc_hd__buf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 1.075000 1.240000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.855000 0.255000 2.025000 0.735000 ;
        RECT 1.855000 0.735000 4.545000 0.905000 ;
        RECT 1.855000 1.445000 4.545000 1.615000 ;
        RECT 1.855000 1.615000 2.025000 2.465000 ;
        RECT 2.695000 0.255000 2.865000 0.735000 ;
        RECT 2.695000 1.615000 2.865000 2.465000 ;
        RECT 3.535000 0.255000 3.705000 0.735000 ;
        RECT 3.535000 1.615000 3.705000 2.465000 ;
        RECT 4.290000 0.905000 4.545000 1.445000 ;
        RECT 4.375000 0.255000 4.545000 0.735000 ;
        RECT 4.375000 1.615000 4.545000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.095000  1.445000 1.595000 1.615000 ;
      RECT 0.095000  1.615000 0.425000 2.465000 ;
      RECT 0.175000  0.255000 0.345000 0.735000 ;
      RECT 0.175000  0.735000 1.595000 0.905000 ;
      RECT 0.515000  0.085000 0.845000 0.565000 ;
      RECT 0.595000  1.835000 0.765000 2.635000 ;
      RECT 0.935000  1.615000 1.265000 2.465000 ;
      RECT 1.015000  0.260000 1.185000 0.735000 ;
      RECT 1.355000  0.085000 1.685000 0.565000 ;
      RECT 1.420000  0.905000 1.595000 1.075000 ;
      RECT 1.420000  1.075000 4.045000 1.245000 ;
      RECT 1.420000  1.245000 1.595000 1.445000 ;
      RECT 1.435000  1.835000 1.605000 2.635000 ;
      RECT 2.195000  0.085000 2.525000 0.565000 ;
      RECT 2.195000  1.835000 2.525000 2.635000 ;
      RECT 3.035000  0.085000 3.365000 0.565000 ;
      RECT 3.035000  1.835000 3.365000 2.635000 ;
      RECT 3.875000  0.085000 4.205000 0.565000 ;
      RECT 3.875000  1.835000 4.205000 2.635000 ;
      RECT 4.715000  0.085000 5.045000 0.885000 ;
      RECT 4.715000  1.485000 5.045000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__buf_8
MACRO sky130_fd_sc_hd__buf_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_12 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 1.075000 1.660000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.673000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.275000 0.255000 2.445000 0.735000 ;
        RECT 2.275000 0.735000 6.645000 0.905000 ;
        RECT 2.275000 1.445000 6.645000 1.615000 ;
        RECT 2.275000 1.615000 2.445000 2.465000 ;
        RECT 3.115000 0.255000 3.285000 0.735000 ;
        RECT 3.115000 1.615000 3.285000 2.465000 ;
        RECT 3.955000 0.255000 4.125000 0.735000 ;
        RECT 3.955000 1.615000 4.125000 2.465000 ;
        RECT 4.710000 0.905000 6.645000 1.445000 ;
        RECT 4.795000 0.255000 4.965000 0.735000 ;
        RECT 4.795000 1.615000 4.965000 2.465000 ;
        RECT 5.635000 0.255000 5.805000 0.735000 ;
        RECT 5.635000 1.615000 5.805000 2.465000 ;
        RECT 6.475000 0.255000 6.645000 0.735000 ;
        RECT 6.475000 1.615000 6.645000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.570000 -0.085000 0.740000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.565000 ;
      RECT 0.175000  1.835000 0.345000 2.635000 ;
      RECT 0.515000  1.445000 2.015000 1.615000 ;
      RECT 0.515000  1.615000 0.845000 2.465000 ;
      RECT 0.595000  0.255000 0.765000 0.735000 ;
      RECT 0.595000  0.735000 2.015000 0.905000 ;
      RECT 0.935000  0.085000 1.265000 0.565000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.355000  1.615000 1.685000 2.465000 ;
      RECT 1.435000  0.260000 1.605000 0.735000 ;
      RECT 1.775000  0.085000 2.105000 0.565000 ;
      RECT 1.840000  0.905000 2.015000 1.075000 ;
      RECT 1.840000  1.075000 4.465000 1.245000 ;
      RECT 1.840000  1.245000 2.015000 1.445000 ;
      RECT 1.855000  1.835000 2.025000 2.635000 ;
      RECT 2.615000  0.085000 2.945000 0.565000 ;
      RECT 2.615000  1.835000 2.945000 2.635000 ;
      RECT 3.455000  0.085000 3.785000 0.565000 ;
      RECT 3.455000  1.835000 3.785000 2.635000 ;
      RECT 4.295000  0.085000 4.625000 0.565000 ;
      RECT 4.295000  1.835000 4.625000 2.635000 ;
      RECT 5.135000  0.085000 5.465000 0.565000 ;
      RECT 5.135000  1.835000 5.465000 2.635000 ;
      RECT 5.975000  0.085000 6.305000 0.565000 ;
      RECT 5.975000  1.835000 6.305000 2.635000 ;
      RECT 6.815000  0.085000 7.145000 0.885000 ;
      RECT 6.815000  1.485000 7.145000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__buf_12
MACRO sky130_fd_sc_hd__buf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.485000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 2.485000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035000 0.255000  3.285000 0.260000 ;
        RECT 3.035000 0.260000  3.365000 0.735000 ;
        RECT 3.035000 0.735000 10.035000 0.905000 ;
        RECT 3.035000 1.445000 10.035000 1.615000 ;
        RECT 3.035000 1.615000  3.365000 2.465000 ;
        RECT 3.875000 0.260000  4.205000 0.735000 ;
        RECT 3.875000 1.615000  4.205000 2.465000 ;
        RECT 3.955000 0.255000  4.125000 0.260000 ;
        RECT 4.715000 0.260000  5.045000 0.735000 ;
        RECT 4.715000 1.615000  5.045000 2.465000 ;
        RECT 4.795000 0.255000  4.965000 0.260000 ;
        RECT 5.555000 0.260000  5.885000 0.735000 ;
        RECT 5.555000 1.615000  5.885000 2.465000 ;
        RECT 6.395000 0.260000  6.725000 0.735000 ;
        RECT 6.395000 1.615000  6.725000 2.465000 ;
        RECT 7.235000 0.260000  7.565000 0.735000 ;
        RECT 7.235000 1.615000  7.565000 2.465000 ;
        RECT 8.075000 0.260000  8.405000 0.735000 ;
        RECT 8.075000 1.615000  8.405000 2.465000 ;
        RECT 8.915000 0.260000  9.245000 0.735000 ;
        RECT 8.915000 1.615000  9.245000 2.465000 ;
        RECT 9.655000 0.905000 10.035000 1.445000 ;
        RECT 9.760000 0.365000 10.035000 0.735000 ;
        RECT 9.760000 1.615000 10.035000 2.360000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.175000  0.085000  0.345000 0.905000 ;
      RECT 0.175000  1.445000  0.345000 2.635000 ;
      RECT 0.515000  0.260000  0.845000 0.735000 ;
      RECT 0.515000  0.735000  2.865000 0.905000 ;
      RECT 0.515000  1.445000  2.865000 1.615000 ;
      RECT 0.515000  1.615000  0.845000 2.465000 ;
      RECT 1.015000  0.085000  1.185000 0.565000 ;
      RECT 1.015000  1.835000  1.185000 2.635000 ;
      RECT 1.355000  0.260000  1.685000 0.735000 ;
      RECT 1.355000  1.615000  1.685000 2.465000 ;
      RECT 1.855000  0.085000  2.025000 0.565000 ;
      RECT 1.855000  1.835000  2.025000 2.635000 ;
      RECT 2.195000  0.260000  2.525000 0.735000 ;
      RECT 2.195000  1.615000  2.525000 2.465000 ;
      RECT 2.690000  0.905000  2.865000 1.075000 ;
      RECT 2.690000  1.075000  9.410000 1.275000 ;
      RECT 2.690000  1.275000  2.865000 1.445000 ;
      RECT 2.695000  0.085000  2.865000 0.565000 ;
      RECT 2.695000  1.835000  2.865000 2.635000 ;
      RECT 3.535000  0.085000  3.705000 0.565000 ;
      RECT 3.535000  1.835000  3.705000 2.635000 ;
      RECT 4.375000  0.085000  4.545000 0.565000 ;
      RECT 4.375000  1.835000  4.545000 2.635000 ;
      RECT 5.215000  0.085000  5.385000 0.565000 ;
      RECT 5.215000  1.835000  5.385000 2.635000 ;
      RECT 6.055000  0.085000  6.225000 0.565000 ;
      RECT 6.055000  1.835000  6.225000 2.635000 ;
      RECT 6.895000  0.085000  7.065000 0.565000 ;
      RECT 6.895000  1.835000  7.065000 2.635000 ;
      RECT 7.735000  0.085000  7.905000 0.565000 ;
      RECT 7.735000  1.835000  7.905000 2.635000 ;
      RECT 8.575000  0.085000  8.745000 0.565000 ;
      RECT 8.575000  1.835000  8.745000 2.635000 ;
      RECT 9.415000  0.085000  9.585000 0.565000 ;
      RECT 9.415000  1.835000  9.585000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
END sky130_fd_sc_hd__buf_16
MACRO sky130_fd_sc_hd__bufbuf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__bufbuf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.230000 0.260000 3.560000 0.735000 ;
        RECT 3.230000 0.735000 6.815000 0.905000 ;
        RECT 3.230000 1.445000 6.815000 1.615000 ;
        RECT 3.230000 1.615000 3.560000 2.465000 ;
        RECT 4.070000 0.260000 4.400000 0.735000 ;
        RECT 4.070000 1.615000 4.400000 2.465000 ;
        RECT 4.910000 0.260000 5.240000 0.735000 ;
        RECT 4.910000 1.615000 5.240000 2.465000 ;
        RECT 5.750000 0.260000 6.080000 0.735000 ;
        RECT 5.750000 1.615000 6.080000 2.465000 ;
        RECT 6.435000 0.905000 6.815000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.090000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.095000  0.260000 0.425000 0.735000 ;
      RECT 0.095000  0.735000 0.780000 0.905000 ;
      RECT 0.095000  1.445000 0.780000 1.615000 ;
      RECT 0.095000  1.615000 0.425000 2.160000 ;
      RECT 0.595000  0.085000 0.765000 0.565000 ;
      RECT 0.595000  1.785000 0.765000 2.635000 ;
      RECT 0.610000  0.905000 0.780000 0.995000 ;
      RECT 0.610000  0.995000 1.040000 1.325000 ;
      RECT 0.610000  1.325000 0.780000 1.445000 ;
      RECT 1.000000  0.260000 1.380000 0.825000 ;
      RECT 1.000000  1.545000 1.380000 2.465000 ;
      RECT 1.210000  0.825000 1.380000 1.075000 ;
      RECT 1.210000  1.075000 2.720000 1.275000 ;
      RECT 1.210000  1.275000 1.380000 1.545000 ;
      RECT 1.550000  0.260000 1.880000 0.735000 ;
      RECT 1.550000  0.735000 3.060000 0.905000 ;
      RECT 1.550000  1.445000 3.060000 1.615000 ;
      RECT 1.550000  1.615000 1.880000 2.465000 ;
      RECT 2.050000  0.085000 2.220000 0.565000 ;
      RECT 2.050000  1.785000 2.220000 2.635000 ;
      RECT 2.390000  0.260000 2.720000 0.735000 ;
      RECT 2.390000  1.615000 2.720000 2.465000 ;
      RECT 2.890000  0.085000 3.060000 0.565000 ;
      RECT 2.890000  0.905000 3.060000 1.075000 ;
      RECT 2.890000  1.075000 5.360000 1.275000 ;
      RECT 2.890000  1.275000 3.060000 1.445000 ;
      RECT 2.890000  1.785000 3.060000 2.635000 ;
      RECT 3.730000  0.085000 3.900000 0.565000 ;
      RECT 3.730000  1.835000 3.900000 2.635000 ;
      RECT 4.570000  0.085000 4.740000 0.565000 ;
      RECT 4.570000  1.835000 4.740000 2.635000 ;
      RECT 5.410000  0.085000 5.580000 0.565000 ;
      RECT 5.410000  1.835000 5.580000 2.635000 ;
      RECT 6.250000  0.085000 6.420000 0.565000 ;
      RECT 6.250000  1.835000 6.420000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
END sky130_fd_sc_hd__bufbuf_8
MACRO sky130_fd_sc_hd__bufbuf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__bufbuf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  5.235000 0.255000  5.485000 0.260000 ;
        RECT  5.235000 0.260000  5.565000 0.735000 ;
        RECT  5.235000 0.735000 11.875000 0.905000 ;
        RECT  5.235000 1.445000 11.875000 1.615000 ;
        RECT  5.235000 1.615000  5.565000 2.465000 ;
        RECT  6.075000 0.260000  6.405000 0.735000 ;
        RECT  6.075000 1.615000  6.405000 2.465000 ;
        RECT  6.155000 0.255000  6.325000 0.260000 ;
        RECT  6.915000 0.260000  7.245000 0.735000 ;
        RECT  6.915000 1.615000  7.245000 2.465000 ;
        RECT  6.995000 0.255000  7.165000 0.260000 ;
        RECT  7.755000 0.260000  8.085000 0.735000 ;
        RECT  7.755000 1.615000  8.085000 2.465000 ;
        RECT  8.595000 0.260000  8.925000 0.735000 ;
        RECT  8.595000 1.615000  8.925000 2.465000 ;
        RECT  9.435000 0.260000  9.765000 0.735000 ;
        RECT  9.435000 1.615000  9.765000 2.465000 ;
        RECT 10.275000 0.260000 10.605000 0.735000 ;
        RECT 10.275000 1.615000 10.605000 2.465000 ;
        RECT 11.115000 0.260000 11.445000 0.735000 ;
        RECT 11.115000 1.615000 11.445000 2.465000 ;
        RECT 11.620000 0.905000 11.875000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.150000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.175000  0.085000  0.345000 0.905000 ;
      RECT  0.175000  1.445000  0.345000 2.635000 ;
      RECT  0.515000  0.260000  0.845000 0.905000 ;
      RECT  0.515000  1.445000  0.845000 2.465000 ;
      RECT  0.610000  0.905000  0.845000 1.075000 ;
      RECT  0.610000  1.075000  2.205000 1.275000 ;
      RECT  0.610000  1.275000  0.845000 1.445000 ;
      RECT  1.035000  0.260000  1.365000 0.735000 ;
      RECT  1.035000  0.735000  2.545000 0.905000 ;
      RECT  1.035000  1.445000  2.545000 1.615000 ;
      RECT  1.035000  1.615000  1.365000 2.465000 ;
      RECT  1.535000  0.085000  1.705000 0.565000 ;
      RECT  1.535000  1.785000  1.705000 2.635000 ;
      RECT  1.875000  0.260000  2.205000 0.735000 ;
      RECT  1.875000  1.615000  2.205000 2.465000 ;
      RECT  2.375000  0.085000  2.545000 0.565000 ;
      RECT  2.375000  0.905000  2.545000 1.075000 ;
      RECT  2.375000  1.075000  4.685000 1.275000 ;
      RECT  2.375000  1.275000  2.545000 1.445000 ;
      RECT  2.375000  1.785000  2.545000 2.635000 ;
      RECT  2.715000  0.260000  3.045000 0.735000 ;
      RECT  2.715000  0.735000  5.065000 0.905000 ;
      RECT  2.715000  1.445000  5.065000 1.615000 ;
      RECT  2.715000  1.615000  3.045000 2.465000 ;
      RECT  3.215000  0.085000  3.385000 0.565000 ;
      RECT  3.215000  1.835000  3.385000 2.635000 ;
      RECT  3.555000  0.260000  3.885000 0.735000 ;
      RECT  3.555000  1.615000  3.885000 2.465000 ;
      RECT  4.055000  0.085000  4.225000 0.565000 ;
      RECT  4.055000  1.835000  4.225000 2.635000 ;
      RECT  4.395000  0.260000  4.725000 0.735000 ;
      RECT  4.395000  1.615000  4.725000 2.465000 ;
      RECT  4.890000  0.905000  5.065000 1.075000 ;
      RECT  4.890000  1.075000 11.450000 1.275000 ;
      RECT  4.890000  1.275000  5.065000 1.445000 ;
      RECT  4.895000  0.085000  5.065000 0.565000 ;
      RECT  4.895000  1.835000  5.065000 2.635000 ;
      RECT  5.735000  0.085000  5.905000 0.565000 ;
      RECT  5.735000  1.835000  5.905000 2.635000 ;
      RECT  6.575000  0.085000  6.745000 0.565000 ;
      RECT  6.575000  1.835000  6.745000 2.635000 ;
      RECT  7.415000  0.085000  7.585000 0.565000 ;
      RECT  7.415000  1.835000  7.585000 2.635000 ;
      RECT  8.255000  0.085000  8.425000 0.565000 ;
      RECT  8.255000  1.835000  8.425000 2.635000 ;
      RECT  9.095000  0.085000  9.265000 0.565000 ;
      RECT  9.095000  1.835000  9.265000 2.635000 ;
      RECT  9.935000  0.085000 10.105000 0.565000 ;
      RECT  9.935000  1.835000 10.105000 2.635000 ;
      RECT 10.775000  0.085000 10.945000 0.565000 ;
      RECT 10.775000  1.835000 10.945000 2.635000 ;
      RECT 11.615000  0.085000 11.785000 0.565000 ;
      RECT 11.615000  1.835000 11.785000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
  END
END sky130_fd_sc_hd__bufbuf_16
MACRO sky130_fd_sc_hd__bufinv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__bufinv_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.505000 1.275000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.715000 0.260000 3.045000 0.735000 ;
        RECT 2.715000 0.735000 6.355000 0.905000 ;
        RECT 2.715000 1.445000 6.355000 1.615000 ;
        RECT 2.715000 1.615000 3.045000 2.465000 ;
        RECT 3.555000 0.260000 3.885000 0.735000 ;
        RECT 3.555000 1.615000 3.885000 2.465000 ;
        RECT 4.395000 0.260000 4.725000 0.735000 ;
        RECT 4.395000 1.615000 4.725000 2.465000 ;
        RECT 5.235000 0.260000 5.565000 0.735000 ;
        RECT 5.235000 1.615000 5.565000 2.465000 ;
        RECT 5.970000 0.905000 6.355000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.175000  0.085000 0.345000 0.905000 ;
      RECT 0.175000  1.445000 0.345000 2.635000 ;
      RECT 0.515000  0.260000 0.845000 0.905000 ;
      RECT 0.515000  1.545000 0.845000 2.465000 ;
      RECT 0.675000  0.905000 0.845000 1.075000 ;
      RECT 0.675000  1.075000 2.205000 1.275000 ;
      RECT 0.675000  1.275000 0.845000 1.545000 ;
      RECT 1.035000  0.260000 1.365000 0.735000 ;
      RECT 1.035000  0.735000 2.545000 0.905000 ;
      RECT 1.035000  1.445000 2.545000 1.615000 ;
      RECT 1.035000  1.615000 1.365000 2.465000 ;
      RECT 1.535000  0.085000 1.705000 0.565000 ;
      RECT 1.535000  1.785000 1.705000 2.635000 ;
      RECT 1.875000  0.260000 2.205000 0.735000 ;
      RECT 1.875000  1.615000 2.205000 2.465000 ;
      RECT 2.375000  0.085000 2.545000 0.565000 ;
      RECT 2.375000  0.905000 2.545000 1.075000 ;
      RECT 2.375000  1.075000 5.760000 1.275000 ;
      RECT 2.375000  1.275000 2.545000 1.445000 ;
      RECT 2.375000  1.785000 2.545000 2.635000 ;
      RECT 3.215000  0.085000 3.385000 0.565000 ;
      RECT 3.215000  1.835000 3.385000 2.635000 ;
      RECT 4.055000  0.085000 4.225000 0.565000 ;
      RECT 4.055000  1.835000 4.225000 2.635000 ;
      RECT 4.895000  0.085000 5.065000 0.565000 ;
      RECT 4.895000  1.835000 5.065000 2.635000 ;
      RECT 5.735000  0.085000 5.905000 0.565000 ;
      RECT 5.735000  1.835000 5.905000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__bufinv_8
MACRO sky130_fd_sc_hd__bufinv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__bufinv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.265000 1.275000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  4.295000 0.255000  4.545000 0.260000 ;
        RECT  4.295000 0.260000  4.625000 0.735000 ;
        RECT  4.295000 0.735000 10.955000 0.905000 ;
        RECT  4.295000 1.445000 10.955000 1.615000 ;
        RECT  4.295000 1.615000  4.625000 2.465000 ;
        RECT  5.135000 0.260000  5.465000 0.735000 ;
        RECT  5.135000 1.615000  5.465000 2.465000 ;
        RECT  5.215000 0.255000  5.385000 0.260000 ;
        RECT  5.975000 0.260000  6.305000 0.735000 ;
        RECT  5.975000 1.615000  6.305000 2.465000 ;
        RECT  6.055000 0.255000  6.225000 0.260000 ;
        RECT  6.815000 0.260000  7.145000 0.735000 ;
        RECT  6.815000 1.615000  7.145000 2.465000 ;
        RECT  7.655000 0.260000  7.985000 0.735000 ;
        RECT  7.655000 1.615000  7.985000 2.465000 ;
        RECT  8.495000 0.260000  8.825000 0.735000 ;
        RECT  8.495000 1.615000  8.825000 2.465000 ;
        RECT  9.335000 0.260000  9.665000 0.735000 ;
        RECT  9.335000 1.615000  9.665000 2.465000 ;
        RECT 10.175000 0.260000 10.505000 0.735000 ;
        RECT 10.175000 1.615000 10.505000 2.465000 ;
        RECT 10.680000 0.905000 10.955000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.095000  0.260000  0.425000 0.735000 ;
      RECT  0.095000  0.735000  1.605000 0.905000 ;
      RECT  0.095000  1.445000  1.605000 1.615000 ;
      RECT  0.095000  1.615000  0.425000 2.465000 ;
      RECT  0.595000  0.085000  0.765000 0.565000 ;
      RECT  0.595000  1.785000  0.765000 2.635000 ;
      RECT  0.935000  0.260000  1.265000 0.735000 ;
      RECT  0.935000  1.615000  1.265000 2.465000 ;
      RECT  1.435000  0.085000  1.605000 0.565000 ;
      RECT  1.435000  0.905000  1.605000 1.075000 ;
      RECT  1.435000  1.075000  3.745000 1.275000 ;
      RECT  1.435000  1.275000  1.605000 1.445000 ;
      RECT  1.435000  1.785000  1.605000 2.635000 ;
      RECT  1.775000  0.260000  2.105000 0.735000 ;
      RECT  1.775000  0.735000  4.125000 0.905000 ;
      RECT  1.775000  1.445000  4.125000 1.615000 ;
      RECT  1.775000  1.615000  2.105000 2.465000 ;
      RECT  2.275000  0.085000  2.445000 0.565000 ;
      RECT  2.275000  1.835000  2.445000 2.635000 ;
      RECT  2.615000  0.260000  2.945000 0.735000 ;
      RECT  2.615000  1.615000  2.945000 2.465000 ;
      RECT  3.115000  0.085000  3.285000 0.565000 ;
      RECT  3.115000  1.835000  3.285000 2.635000 ;
      RECT  3.455000  0.260000  3.785000 0.735000 ;
      RECT  3.455000  1.615000  3.785000 2.465000 ;
      RECT  3.950000  0.905000  4.125000 1.075000 ;
      RECT  3.950000  1.075000 10.510000 1.275000 ;
      RECT  3.950000  1.275000  4.125000 1.445000 ;
      RECT  3.955000  0.085000  4.125000 0.565000 ;
      RECT  3.955000  1.835000  4.125000 2.635000 ;
      RECT  4.795000  0.085000  4.965000 0.565000 ;
      RECT  4.795000  1.835000  4.965000 2.635000 ;
      RECT  5.635000  0.085000  5.805000 0.565000 ;
      RECT  5.635000  1.835000  5.805000 2.635000 ;
      RECT  6.475000  0.085000  6.645000 0.565000 ;
      RECT  6.475000  1.835000  6.645000 2.635000 ;
      RECT  7.315000  0.085000  7.485000 0.565000 ;
      RECT  7.315000  1.835000  7.485000 2.635000 ;
      RECT  8.155000  0.085000  8.325000 0.565000 ;
      RECT  8.155000  1.835000  8.325000 2.635000 ;
      RECT  8.995000  0.085000  9.165000 0.565000 ;
      RECT  8.995000  1.835000  9.165000 2.635000 ;
      RECT  9.835000  0.085000 10.005000 0.565000 ;
      RECT  9.835000  1.835000 10.005000 2.635000 ;
      RECT 10.675000  0.085000 10.845000 0.565000 ;
      RECT 10.675000  1.835000 10.845000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
  END
END sky130_fd_sc_hd__bufinv_16
MACRO sky130_fd_sc_hd__clkbuf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.196500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.985000 1.275000 1.355000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.345000 0.760000 ;
        RECT 0.085000 0.760000 0.255000 1.560000 ;
        RECT 0.085000 1.560000 0.355000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.425000  1.060000 0.710000 1.390000 ;
      RECT 0.525000  0.085000 0.855000 0.465000 ;
      RECT 0.525000  1.875000 0.855000 2.635000 ;
      RECT 0.540000  0.635000 1.205000 0.805000 ;
      RECT 0.540000  0.805000 0.710000 1.060000 ;
      RECT 0.540000  1.390000 0.710000 1.535000 ;
      RECT 0.540000  1.535000 1.205000 1.705000 ;
      RECT 1.035000  0.255000 1.205000 0.635000 ;
      RECT 1.035000  1.705000 1.205000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__clkbuf_1
MACRO sky130_fd_sc_hd__clkbuf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.745000 0.785000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.383400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.040000 0.255000 1.245000 0.655000 ;
        RECT 1.040000 0.655000 1.725000 0.825000 ;
        RECT 1.060000 1.855000 1.725000 2.030000 ;
        RECT 1.060000 2.030000 1.245000 2.435000 ;
        RECT 1.385000 0.825000 1.725000 1.855000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.585000 ;
      RECT 0.085000  0.585000 0.255000 1.495000 ;
      RECT 0.085000  1.495000 1.215000 1.665000 ;
      RECT 0.085000  1.665000 0.355000 2.435000 ;
      RECT 0.525000  1.855000 0.855000 2.635000 ;
      RECT 0.555000  0.085000 0.830000 0.565000 ;
      RECT 0.965000  0.995000 1.215000 1.495000 ;
      RECT 1.415000  0.085000 1.750000 0.485000 ;
      RECT 1.415000  2.210000 1.750000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__clkbuf_2
MACRO sky130_fd_sc_hd__clkbuf_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.755000 0.775000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.795200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.345000 1.305000 0.735000 ;
        RECT 1.010000 0.735000 2.660000 0.905000 ;
        RECT 1.045000 1.835000 2.165000 2.005000 ;
        RECT 1.045000 2.005000 1.305000 2.465000 ;
        RECT 1.905000 0.345000 2.165000 0.735000 ;
        RECT 1.905000 1.415000 2.660000 1.585000 ;
        RECT 1.905000 1.585000 2.165000 1.835000 ;
        RECT 1.905000 2.005000 2.165000 2.465000 ;
        RECT 2.255000 0.905000 2.660000 1.415000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.255000 0.385000 0.585000 ;
      RECT 0.085000  0.585000 0.255000 1.495000 ;
      RECT 0.085000  1.495000 1.115000 1.665000 ;
      RECT 0.085000  1.665000 0.395000 2.465000 ;
      RECT 0.555000  0.085000 0.830000 0.565000 ;
      RECT 0.565000  1.835000 0.875000 2.635000 ;
      RECT 0.945000  1.075000 2.085000 1.245000 ;
      RECT 0.945000  1.245000 1.115000 1.495000 ;
      RECT 1.475000  0.085000 1.730000 0.565000 ;
      RECT 1.475000  2.175000 1.730000 2.635000 ;
      RECT 2.335000  0.085000 2.615000 0.565000 ;
      RECT 2.335000  1.765000 2.620000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__clkbuf_4
MACRO sky130_fd_sc_hd__clkbuf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.426000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 0.400000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.590400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.420000 0.280000 1.680000 0.735000 ;
        RECT 1.420000 0.735000 4.730000 0.905000 ;
        RECT 1.420000 1.495000 4.730000 1.735000 ;
        RECT 1.420000 1.735000 1.680000 2.460000 ;
        RECT 2.280000 0.280000 2.540000 0.735000 ;
        RECT 2.280000 1.735000 2.540000 2.460000 ;
        RECT 3.140000 0.280000 3.400000 0.735000 ;
        RECT 3.140000 1.735000 3.400000 2.460000 ;
        RECT 3.760000 0.905000 4.730000 1.495000 ;
        RECT 4.000000 0.280000 4.260000 0.735000 ;
        RECT 4.000000 1.735000 4.260000 2.460000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.095000  1.525000 0.390000 2.635000 ;
      RECT 0.145000  0.085000 0.390000 0.545000 ;
      RECT 0.570000  0.265000 0.820000 1.075000 ;
      RECT 0.570000  1.075000 3.590000 1.325000 ;
      RECT 0.570000  1.325000 0.820000 2.460000 ;
      RECT 0.990000  0.085000 1.250000 0.610000 ;
      RECT 0.990000  1.525000 1.250000 2.635000 ;
      RECT 1.850000  0.085000 2.110000 0.565000 ;
      RECT 1.850000  1.905000 2.110000 2.635000 ;
      RECT 2.710000  0.085000 2.970000 0.565000 ;
      RECT 2.710000  1.905000 2.970000 2.635000 ;
      RECT 3.570000  0.085000 3.830000 0.565000 ;
      RECT 3.570000  1.905000 3.830000 2.635000 ;
      RECT 4.430000  0.085000 4.730000 0.565000 ;
      RECT 4.430000  1.905000 4.725000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__clkbuf_8
MACRO sky130_fd_sc_hd__clkbuf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.852000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.400000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.180800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.280000 0.280000 2.540000 0.735000 ;
        RECT 2.280000 0.735000 9.025000 0.905000 ;
        RECT 2.280000 1.495000 9.025000 1.720000 ;
        RECT 2.280000 1.720000 7.685000 1.735000 ;
        RECT 2.280000 1.735000 2.540000 2.460000 ;
        RECT 3.140000 0.280000 3.400000 0.735000 ;
        RECT 3.140000 1.735000 3.400000 2.460000 ;
        RECT 4.000000 0.280000 4.260000 0.735000 ;
        RECT 4.000000 1.735000 4.260000 2.460000 ;
        RECT 4.845000 0.280000 5.120000 0.735000 ;
        RECT 4.860000 1.735000 5.120000 2.460000 ;
        RECT 5.705000 0.280000 5.965000 0.735000 ;
        RECT 5.705000 1.735000 5.965000 2.460000 ;
        RECT 6.565000 0.280000 6.825000 0.735000 ;
        RECT 6.565000 1.735000 6.825000 2.460000 ;
        RECT 7.425000 0.280000 7.685000 0.735000 ;
        RECT 7.425000 1.735000 7.685000 2.460000 ;
        RECT 7.860000 0.905000 9.025000 1.495000 ;
        RECT 8.295000 0.280000 8.555000 0.735000 ;
        RECT 8.295000 1.720000 8.585000 2.460000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.085000  0.085000 0.390000 0.595000 ;
      RECT 0.095000  1.825000 0.390000 2.635000 ;
      RECT 0.570000  0.265000 0.820000 1.075000 ;
      RECT 0.570000  1.075000 7.690000 1.325000 ;
      RECT 0.570000  1.325000 0.815000 2.465000 ;
      RECT 0.990000  0.085000 1.250000 0.610000 ;
      RECT 0.990000  1.825000 1.250000 2.635000 ;
      RECT 1.430000  0.265000 1.680000 1.075000 ;
      RECT 1.430000  1.325000 1.680000 2.460000 ;
      RECT 1.850000  0.085000 2.110000 0.645000 ;
      RECT 1.850000  1.835000 2.110000 2.630000 ;
      RECT 1.850000  2.630000 8.125000 2.635000 ;
      RECT 2.710000  0.085000 2.970000 0.565000 ;
      RECT 2.710000  1.905000 2.970000 2.630000 ;
      RECT 3.570000  0.085000 3.830000 0.565000 ;
      RECT 3.570000  1.905000 3.830000 2.630000 ;
      RECT 4.430000  0.085000 4.675000 0.565000 ;
      RECT 4.430000  1.905000 4.690000 2.630000 ;
      RECT 5.290000  0.085000 5.535000 0.565000 ;
      RECT 5.290000  1.905000 5.535000 2.630000 ;
      RECT 6.145000  0.085000 6.395000 0.565000 ;
      RECT 6.150000  1.905000 6.395000 2.630000 ;
      RECT 7.005000  0.085000 7.255000 0.565000 ;
      RECT 7.010000  1.905000 7.255000 2.630000 ;
      RECT 7.865000  0.085000 8.125000 0.565000 ;
      RECT 7.870000  1.905000 8.125000 2.630000 ;
      RECT 8.725000  0.085000 9.025000 0.565000 ;
      RECT 8.755000  1.890000 9.025000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
  END
END sky130_fd_sc_hd__clkbuf_16
MACRO sky130_fd_sc_hd__clkdlybuf4s15_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s15_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.560000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.376300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.210000 0.285000 3.595000 0.545000 ;
        RECT 3.210000 1.760000 3.595000 2.465000 ;
        RECT 3.365000 0.545000 3.595000 1.760000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.255000 0.425000 0.715000 ;
      RECT 0.085000  0.715000 1.215000 0.885000 ;
      RECT 0.085000  1.495000 1.215000 1.665000 ;
      RECT 0.085000  1.665000 0.425000 2.465000 ;
      RECT 0.595000  0.085000 0.910000 0.545000 ;
      RECT 0.595000  1.835000 0.925000 2.635000 ;
      RECT 0.730000  0.885000 1.215000 1.495000 ;
      RECT 1.385000  0.255000 1.760000 0.825000 ;
      RECT 1.385000  1.835000 1.760000 2.465000 ;
      RECT 1.590000  0.825000 1.760000 1.055000 ;
      RECT 1.590000  1.055000 2.685000 1.250000 ;
      RECT 1.590000  1.250000 1.760000 1.835000 ;
      RECT 1.930000  0.255000 2.260000 0.715000 ;
      RECT 1.930000  0.715000 3.195000 0.885000 ;
      RECT 1.930000  1.420000 3.195000 1.590000 ;
      RECT 1.930000  1.590000 2.410000 2.465000 ;
      RECT 2.640000  1.760000 3.040000 2.635000 ;
      RECT 2.710000  0.085000 3.040000 0.545000 ;
      RECT 2.855000  0.885000 3.195000 1.420000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s15_1
MACRO sky130_fd_sc_hd__clkdlybuf4s15_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s15_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.060000 0.555000 1.625000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.397600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.050000 0.255000 3.550000 0.640000 ;
        RECT 3.070000 1.485000 3.550000 2.465000 ;
        RECT 3.355000 0.640000 3.550000 1.485000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.255000 0.415000 0.720000 ;
      RECT 0.085000  0.720000 1.060000 0.890000 ;
      RECT 0.085000  1.795000 1.060000 1.965000 ;
      RECT 0.085000  1.965000 0.430000 2.465000 ;
      RECT 0.585000  0.085000 0.915000 0.550000 ;
      RECT 0.600000  2.135000 0.930000 2.635000 ;
      RECT 0.890000  0.890000 1.060000 1.075000 ;
      RECT 0.890000  1.075000 1.320000 1.245000 ;
      RECT 0.890000  1.245000 1.060000 1.795000 ;
      RECT 1.230000  1.785000 1.660000 2.465000 ;
      RECT 1.280000  0.255000 1.660000 0.905000 ;
      RECT 1.490000  0.905000 1.660000 1.075000 ;
      RECT 1.490000  1.075000 2.415000 1.485000 ;
      RECT 1.490000  1.485000 1.660000 1.785000 ;
      RECT 1.830000  0.255000 2.100000 0.735000 ;
      RECT 1.830000  0.735000 2.900000 0.905000 ;
      RECT 1.830000  1.790000 2.900000 1.965000 ;
      RECT 1.830000  1.965000 2.100000 2.465000 ;
      RECT 2.550000  0.085000 2.880000 0.565000 ;
      RECT 2.550000  2.135000 2.880000 2.635000 ;
      RECT 2.730000  0.905000 2.900000 1.075000 ;
      RECT 2.730000  1.075000 3.185000 1.245000 ;
      RECT 2.730000  1.245000 2.900000 1.790000 ;
      RECT 3.720000  0.085000 4.055000 0.645000 ;
      RECT 3.720000  1.485000 4.055000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s15_2
MACRO sky130_fd_sc_hd__clkdlybuf4s18_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s18_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.055000 0.550000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.376300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.210000 0.255000 3.590000 0.545000 ;
        RECT 3.220000 1.760000 3.590000 2.465000 ;
        RECT 3.365000 0.545000 3.590000 1.760000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.095000  0.255000 0.425000 0.715000 ;
      RECT 0.095000  0.715000 1.215000 0.885000 ;
      RECT 0.095000  1.495000 1.215000 1.665000 ;
      RECT 0.095000  1.665000 0.425000 2.465000 ;
      RECT 0.595000  0.085000 0.910000 0.545000 ;
      RECT 0.595000  1.835000 0.925000 2.635000 ;
      RECT 0.720000  0.885000 1.215000 1.495000 ;
      RECT 1.385000  0.255000 1.760000 0.825000 ;
      RECT 1.385000  1.835000 1.760000 2.465000 ;
      RECT 1.590000  0.825000 1.760000 1.055000 ;
      RECT 1.590000  1.055000 2.685000 1.250000 ;
      RECT 1.590000  1.250000 1.760000 1.835000 ;
      RECT 1.930000  0.255000 2.260000 0.715000 ;
      RECT 1.930000  0.715000 3.195000 0.885000 ;
      RECT 1.930000  1.420000 3.195000 1.590000 ;
      RECT 1.930000  1.590000 2.260000 2.465000 ;
      RECT 2.710000  0.085000 3.040000 0.545000 ;
      RECT 2.710000  1.760000 3.040000 2.635000 ;
      RECT 2.855000  0.885000 3.195000 1.420000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s18_1
MACRO sky130_fd_sc_hd__clkdlybuf4s18_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s18_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.560000 1.290000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.397600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.705000 0.270000 3.150000 0.640000 ;
        RECT 2.715000 1.420000 3.180000 1.525000 ;
        RECT 2.715000 1.525000 3.150000 2.465000 ;
        RECT 2.965000 0.640000 3.150000 0.780000 ;
        RECT 2.965000 0.780000 3.180000 0.945000 ;
        RECT 3.010000 0.945000 3.180000 1.420000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.270000 0.415000 0.735000 ;
      RECT 0.085000  0.735000 1.055000 0.905000 ;
      RECT 0.085000  1.460000 1.055000 1.630000 ;
      RECT 0.085000  1.630000 0.430000 2.465000 ;
      RECT 0.585000  0.085000 0.915000 0.565000 ;
      RECT 0.600000  1.800000 0.930000 2.635000 ;
      RECT 0.730000  0.905000 1.055000 1.460000 ;
      RECT 1.110000  1.800000 1.440000 2.465000 ;
      RECT 1.160000  0.270000 1.440000 0.600000 ;
      RECT 1.270000  0.600000 1.440000 1.075000 ;
      RECT 1.270000  1.075000 2.205000 1.255000 ;
      RECT 1.270000  1.255000 1.440000 1.800000 ;
      RECT 1.630000  0.270000 1.960000 0.735000 ;
      RECT 1.630000  0.735000 2.545000 0.905000 ;
      RECT 1.630000  1.460000 2.545000 1.630000 ;
      RECT 1.630000  1.630000 1.960000 2.465000 ;
      RECT 2.130000  1.800000 2.545000 2.635000 ;
      RECT 2.165000  0.085000 2.535000 0.565000 ;
      RECT 2.375000  0.905000 2.545000 1.075000 ;
      RECT 2.375000  1.075000 2.840000 1.245000 ;
      RECT 2.375000  1.245000 2.545000 1.460000 ;
      RECT 3.320000  0.085000 3.595000 0.645000 ;
      RECT 3.320000  1.625000 3.595000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s18_2
MACRO sky130_fd_sc_hd__clkdlybuf4s25_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s25_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.485000 1.320000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.702900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.015000 0.255000 3.595000 0.640000 ;
        RECT 3.035000 1.565000 3.595000 2.465000 ;
        RECT 3.230000 0.640000 3.595000 1.565000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.255000 0.410000 0.735000 ;
      RECT 0.085000  0.735000 1.005000 0.905000 ;
      RECT 0.085000  1.490000 1.005000 1.660000 ;
      RECT 0.085000  1.660000 0.430000 2.465000 ;
      RECT 0.580000  0.085000 0.910000 0.565000 ;
      RECT 0.600000  1.830000 0.925000 2.635000 ;
      RECT 0.655000  0.905000 1.005000 1.025000 ;
      RECT 0.655000  1.025000 1.105000 1.295000 ;
      RECT 0.655000  1.295000 1.005000 1.490000 ;
      RECT 1.175000  0.255000 1.645000 0.855000 ;
      RECT 1.195000  1.790000 1.645000 2.465000 ;
      RECT 1.470000  0.855000 1.645000 1.075000 ;
      RECT 1.470000  1.075000 2.420000 1.250000 ;
      RECT 1.470000  1.250000 1.645000 1.790000 ;
      RECT 1.815000  0.255000 2.065000 0.735000 ;
      RECT 1.815000  0.735000 2.765000 0.905000 ;
      RECT 1.815000  1.495000 2.765000 1.665000 ;
      RECT 1.815000  1.665000 2.065000 2.465000 ;
      RECT 2.235000  1.835000 2.845000 2.635000 ;
      RECT 2.240000  0.085000 2.845000 0.565000 ;
      RECT 2.595000  0.905000 2.765000 0.990000 ;
      RECT 2.595000  0.990000 3.050000 1.325000 ;
      RECT 2.595000  1.325000 2.765000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s25_1
MACRO sky130_fd_sc_hd__clkdlybuf4s25_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s25_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.495000 1.615000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.497000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.770000 0.285000 3.095000 0.615000 ;
        RECT 2.770000 1.625000 3.095000 2.460000 ;
        RECT 2.865000 0.615000 3.095000 0.765000 ;
        RECT 2.865000 0.765000 3.595000 1.275000 ;
        RECT 2.865000 1.275000 3.095000 1.625000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.095000  0.305000 0.345000 0.640000 ;
      RECT 0.095000  0.640000 0.840000 0.810000 ;
      RECT 0.095000  1.785000 0.835000 1.955000 ;
      RECT 0.095000  1.955000 0.345000 2.465000 ;
      RECT 0.575000  0.085000 0.905000 0.470000 ;
      RECT 0.575000  2.125000 0.905000 2.635000 ;
      RECT 0.665000  0.810000 0.840000 0.995000 ;
      RECT 0.665000  0.995000 1.035000 1.325000 ;
      RECT 0.665000  1.325000 1.005000 1.750000 ;
      RECT 0.665000  1.750000 0.835000 1.785000 ;
      RECT 1.095000  0.255000 1.425000 0.780000 ;
      RECT 1.175000  1.425000 1.440000 2.465000 ;
      RECT 1.205000  0.780000 1.425000 0.995000 ;
      RECT 1.205000  0.995000 2.165000 1.325000 ;
      RECT 1.205000  1.325000 1.440000 1.425000 ;
      RECT 1.615000  0.255000 1.945000 0.635000 ;
      RECT 1.615000  0.635000 2.595000 0.805000 ;
      RECT 1.695000  1.500000 2.595000 1.745000 ;
      RECT 1.695000  1.745000 1.945000 2.465000 ;
      RECT 2.135000  0.085000 2.465000 0.465000 ;
      RECT 2.135000  1.915000 2.465000 2.635000 ;
      RECT 2.335000  0.805000 2.595000 1.500000 ;
      RECT 3.265000  0.085000 3.595000 0.550000 ;
      RECT 3.265000  1.635000 3.595000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s25_2
MACRO sky130_fd_sc_hd__clkdlybuf4s50_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s50_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.535000 1.290000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.190000 0.255000 3.595000 0.640000 ;
        RECT 3.190000 1.690000 3.595000 2.465000 ;
        RECT 3.345000 0.640000 3.595000 1.690000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.255000 0.415000 0.735000 ;
      RECT 0.085000  0.735000 1.055000 0.905000 ;
      RECT 0.085000  1.460000 1.055000 1.630000 ;
      RECT 0.085000  1.630000 0.430000 2.465000 ;
      RECT 0.585000  0.085000 0.915000 0.565000 ;
      RECT 0.600000  1.800000 0.930000 2.635000 ;
      RECT 0.705000  0.905000 1.055000 1.025000 ;
      RECT 0.705000  1.025000 1.135000 1.315000 ;
      RECT 0.705000  1.315000 1.055000 1.460000 ;
      RECT 1.380000  0.255000 1.730000 1.070000 ;
      RECT 1.380000  1.070000 2.240000 1.320000 ;
      RECT 1.380000  1.320000 1.730000 2.465000 ;
      RECT 1.990000  0.255000 2.240000 0.730000 ;
      RECT 1.990000  0.730000 2.580000 0.900000 ;
      RECT 1.990000  1.495000 2.580000 1.665000 ;
      RECT 1.990000  1.665000 2.240000 2.465000 ;
      RECT 2.410000  0.900000 2.580000 0.995000 ;
      RECT 2.410000  0.995000 3.175000 1.325000 ;
      RECT 2.410000  1.325000 2.580000 1.495000 ;
      RECT 2.690000  0.085000 3.020000 0.600000 ;
      RECT 2.690000  1.835000 3.020000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s50_1
MACRO sky130_fd_sc_hd__clkdlybuf4s50_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s50_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.480000 1.285000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.390500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.185000 0.270000 3.625000 0.640000 ;
        RECT 3.185000 1.530000 3.625000 2.465000 ;
        RECT 3.345000 0.640000 3.625000 1.530000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.270000 0.415000 0.735000 ;
      RECT 0.085000  0.735000 1.270000 0.905000 ;
      RECT 0.085000  1.455000 1.270000 1.630000 ;
      RECT 0.085000  1.630000 0.430000 2.465000 ;
      RECT 0.585000  0.085000 0.915000 0.565000 ;
      RECT 0.600000  1.800000 0.930000 2.635000 ;
      RECT 0.765000  1.075000 1.435000 1.245000 ;
      RECT 0.850000  0.905000 1.270000 1.075000 ;
      RECT 0.850000  1.245000 1.270000 1.455000 ;
      RECT 1.390000  1.785000 1.795000 2.465000 ;
      RECT 1.440000  0.270000 1.795000 0.900000 ;
      RECT 1.625000  0.900000 1.795000 1.075000 ;
      RECT 1.625000  1.075000 2.305000 1.245000 ;
      RECT 1.625000  1.245000 1.795000 1.785000 ;
      RECT 1.985000  0.270000 2.235000 0.735000 ;
      RECT 1.985000  0.735000 2.645000 0.905000 ;
      RECT 1.985000  1.460000 2.645000 1.630000 ;
      RECT 1.985000  1.630000 2.235000 2.465000 ;
      RECT 2.475000  0.905000 2.645000 0.995000 ;
      RECT 2.475000  0.995000 3.175000 1.325000 ;
      RECT 2.475000  1.325000 2.645000 1.460000 ;
      RECT 2.685000  0.085000 3.015000 0.565000 ;
      RECT 2.685000  1.800000 3.015000 2.635000 ;
      RECT 3.795000  0.085000 4.055000 0.635000 ;
      RECT 3.795000  1.800000 4.055000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s50_2
MACRO sky130_fd_sc_hd__clkinv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.375000 0.325000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.336000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.840000 0.760000 ;
        RECT 0.515000 0.760000 1.295000 1.290000 ;
        RECT 0.515000 1.290000 0.845000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.085000  1.665000 0.345000 2.635000 ;
      RECT 1.010000  0.085000 1.295000 0.590000 ;
      RECT 1.015000  1.665000 1.295000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__clkinv_1
MACRO sky130_fd_sc_hd__clkinv_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.576000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.065000 1.305000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.662600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.460000 1.755000 1.630000 ;
        RECT 0.155000 1.630000 0.410000 2.435000 ;
        RECT 1.010000 1.630000 1.270000 2.435000 ;
        RECT 1.025000 0.280000 1.250000 0.725000 ;
        RECT 1.025000 0.725000 1.755000 0.895000 ;
        RECT 1.475000 0.895000 1.755000 1.460000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.560000  0.085000 0.855000 0.610000 ;
      RECT 0.580000  1.800000 0.840000 2.635000 ;
      RECT 1.420000  0.085000 1.750000 0.555000 ;
      RECT 1.440000  1.800000 1.695000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__clkinv_2
MACRO sky130_fd_sc_hd__clkinv_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.152000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.065000 2.660000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.075200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.725000 3.135000 0.895000 ;
        RECT 0.105000 0.895000 0.275000 1.460000 ;
        RECT 0.105000 1.460000 3.135000 1.630000 ;
        RECT 0.605000 1.630000 0.860000 2.435000 ;
        RECT 1.030000 0.280000 1.290000 0.725000 ;
        RECT 1.465000 1.630000 1.720000 2.435000 ;
        RECT 1.890000 0.280000 2.145000 0.725000 ;
        RECT 2.320000 1.630000 2.580000 2.435000 ;
        RECT 2.835000 0.895000 3.135000 1.460000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  1.800000 0.430000 2.635000 ;
      RECT 0.565000  0.085000 0.860000 0.555000 ;
      RECT 1.030000  1.800000 1.290000 2.635000 ;
      RECT 1.460000  0.085000 1.720000 0.555000 ;
      RECT 1.890000  1.800000 2.150000 2.635000 ;
      RECT 2.315000  0.085000 2.615000 0.555000 ;
      RECT 2.750000  1.800000 3.135000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__clkinv_4
MACRO sky130_fd_sc_hd__clkinv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.304000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.035000 4.865000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.090400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.695000 5.440000 0.865000 ;
        RECT 0.115000 0.865000 0.285000 1.460000 ;
        RECT 0.115000 1.460000 5.440000 1.630000 ;
        RECT 0.565000 1.630000 0.805000 2.435000 ;
        RECT 1.405000 1.630000 1.645000 2.435000 ;
        RECT 1.535000 0.280000 1.725000 0.695000 ;
        RECT 2.245000 1.630000 2.495000 2.435000 ;
        RECT 2.395000 0.280000 2.585000 0.695000 ;
        RECT 3.080000 1.630000 3.325000 2.435000 ;
        RECT 3.255000 0.280000 3.445000 0.695000 ;
        RECT 3.920000 1.630000 4.175000 2.435000 ;
        RECT 4.115000 0.280000 4.305000 0.695000 ;
        RECT 4.765000 1.630000 5.005000 2.435000 ;
        RECT 5.170000 0.865000 5.440000 1.460000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.135000  1.800000 0.395000 2.635000 ;
      RECT 0.975000  1.800000 1.235000 2.635000 ;
      RECT 1.035000  0.085000 1.365000 0.525000 ;
      RECT 1.815000  1.800000 2.075000 2.635000 ;
      RECT 1.895000  0.085000 2.225000 0.525000 ;
      RECT 2.665000  1.800000 2.910000 2.635000 ;
      RECT 2.755000  0.085000 3.085000 0.525000 ;
      RECT 3.495000  1.800000 3.750000 2.635000 ;
      RECT 3.615000  0.085000 3.945000 0.525000 ;
      RECT 4.345000  1.800000 4.595000 2.635000 ;
      RECT 4.475000  0.085000 4.805000 0.525000 ;
      RECT 5.175000  1.800000 5.430000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__clkinv_8
MACRO sky130_fd_sc_hd__clkinv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  4.608000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.345000 0.895000  2.155000 1.275000 ;
        RECT 8.930000 0.895000 10.710000 1.275000 ;
      LAYER mcon ;
        RECT 1.525000 1.105000 1.695000 1.275000 ;
        RECT 1.985000 1.105000 2.155000 1.275000 ;
        RECT 9.345000 1.105000 9.515000 1.275000 ;
        RECT 9.805000 1.105000 9.975000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465000 1.075000  2.215000 1.120000 ;
        RECT 1.465000 1.120000 10.035000 1.260000 ;
        RECT 1.465000 1.260000  2.215000 1.305000 ;
        RECT 9.285000 1.075000 10.035000 1.120000 ;
        RECT 9.285000 1.260000 10.035000 1.305000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  4.520900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.575000 1.455000 10.480000 1.665000 ;
        RECT  0.575000 1.665000  0.830000 2.465000 ;
        RECT  1.435000 1.665000  1.690000 2.450000 ;
        RECT  2.325000 0.280000  2.550000 1.415000 ;
        RECT  2.325000 1.415000  8.755000 1.455000 ;
        RECT  2.325000 1.665000  2.550000 2.465000 ;
        RECT  3.155000 0.280000  3.410000 1.415000 ;
        RECT  3.155000 1.665000  3.410000 2.450000 ;
        RECT  4.015000 0.280000  4.255000 1.415000 ;
        RECT  4.015000 1.665000  4.255000 2.450000 ;
        RECT  4.905000 0.280000  5.255000 1.415000 ;
        RECT  4.905000 1.665000  5.280000 2.450000 ;
        RECT  5.925000 0.280000  6.175000 1.415000 ;
        RECT  5.925000 1.665000  6.175000 2.450000 ;
        RECT  6.785000 0.280000  7.035000 1.415000 ;
        RECT  6.785000 1.665000  7.035000 2.450000 ;
        RECT  7.645000 0.280000  7.895000 1.415000 ;
        RECT  7.645000 1.665000  7.895000 2.450000 ;
        RECT  8.505000 0.280000  8.755000 1.415000 ;
        RECT  8.505000 1.665000  8.755000 2.450000 ;
        RECT  9.365000 1.665000  9.605000 2.450000 ;
        RECT 10.225000 1.665000 10.480000 2.450000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.140000  1.495000  0.405000 2.635000 ;
      RECT  1.000000  1.835000  1.260000 2.635000 ;
      RECT  1.855000  0.085000  2.125000 0.610000 ;
      RECT  1.865000  1.835000  2.120000 2.635000 ;
      RECT  2.720000  0.085000  2.985000 0.610000 ;
      RECT  2.720000  1.835000  2.980000 2.635000 ;
      RECT  3.580000  0.085000  3.845000 0.610000 ;
      RECT  3.585000  1.835000  3.840000 2.635000 ;
      RECT  4.465000  0.085000  4.730000 0.610000 ;
      RECT  4.465000  1.835000  4.720000 2.635000 ;
      RECT  5.490000  0.085000  5.755000 0.610000 ;
      RECT  5.490000  1.835000  5.745000 2.120000 ;
      RECT  5.490000  2.120000  5.750000 2.635000 ;
      RECT  6.350000  0.085000  6.575000 0.610000 ;
      RECT  6.355000  1.835000  6.610000 2.635000 ;
      RECT  7.210000  0.085000  7.475000 0.610000 ;
      RECT  7.215000  1.835000  7.470000 2.635000 ;
      RECT  8.070000  0.085000  8.335000 0.610000 ;
      RECT  8.075000  1.835000  8.330000 2.635000 ;
      RECT  8.930000  0.085000  9.195000 0.610000 ;
      RECT  8.935000  1.835000  9.190000 2.635000 ;
      RECT  9.795000  1.835000 10.050000 2.635000 ;
      RECT 10.650000  1.835000 10.910000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
  END
END sky130_fd_sc_hd__clkinv_16
MACRO sky130_fd_sc_hd__clkinvlp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinvlp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.995000 0.600000 1.665000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.436750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.810000 0.315000 1.445000 0.750000 ;
        RECT 0.810000 0.750000 1.235000 2.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.225000  1.835000 0.555000 2.625000 ;
      RECT 0.225000  2.625000 1.740000 2.635000 ;
      RECT 0.295000  0.085000 0.625000 0.745000 ;
      RECT 1.440000  1.455000 1.740000 2.625000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__clkinvlp_2
MACRO sky130_fd_sc_hd__clkinvlp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinvlp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.330000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.745000 0.425000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.714000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.255000 1.215000 0.680000 ;
        RECT 0.595000 0.680000 0.955000 1.015000 ;
        RECT 0.595000 1.015000 2.015000 1.295000 ;
        RECT 0.595000 1.295000 0.955000 2.465000 ;
        RECT 1.685000 1.295000 2.015000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.575000 ;
      RECT 0.095000  1.495000 0.425000 2.635000 ;
      RECT 1.155000  1.465000 1.485000 2.635000 ;
      RECT 1.675000  0.085000 2.005000 0.775000 ;
      RECT 2.215000  1.465000 2.545000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__clkinvlp_4
MACRO sky130_fd_sc_hd__conb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__conb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.605000 1.740000 ;
    END
  END HI
  PIN LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.775000 0.915000 1.295000 2.465000 ;
    END
  END LO
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.275000  1.910000 0.605000 2.635000 ;
      RECT 0.775000  0.085000 1.115000 0.745000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__conb_1
MACRO sky130_fd_sc_hd__decap_3
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__decap_3 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.085000  0.085000 1.295000 0.835000 ;
      RECT 0.085000  0.835000 0.605000 1.375000 ;
      RECT 0.085000  1.545000 1.295000 2.635000 ;
      RECT 0.775000  1.005000 1.295000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__decap_3
MACRO sky130_fd_sc_hd__decap_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__decap_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.085000  0.085000 1.755000 0.855000 ;
      RECT 0.085000  0.855000 0.835000 1.375000 ;
      RECT 0.085000  1.545000 1.755000 2.635000 ;
      RECT 1.005000  1.025000 1.755000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__decap_4
MACRO sky130_fd_sc_hd__decap_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__decap_6 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.085000 2.675000 0.855000 ;
      RECT 0.085000  0.855000 1.295000 1.375000 ;
      RECT 0.085000  1.545000 2.675000 2.635000 ;
      RECT 1.465000  1.025000 2.675000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__decap_6
MACRO sky130_fd_sc_hd__decap_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__decap_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.085000 3.595000 0.855000 ;
      RECT 0.085000  0.855000 1.735000 1.375000 ;
      RECT 0.085000  1.545000 3.595000 2.635000 ;
      RECT 1.905000  1.025000 3.595000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__decap_8
MACRO sky130_fd_sc_hd__decap_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__decap_12 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.085000 5.430000 0.855000 ;
      RECT 0.085000  0.855000 2.665000 1.375000 ;
      RECT 0.085000  1.545000 5.430000 2.635000 ;
      RECT 2.835000  1.025000 5.430000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__decap_12
MACRO sky130_fd_sc_hd__dfbbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfbbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.745000 1.005000 2.155000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.615000 0.255000 11.875000 0.825000 ;
        RECT 11.615000 1.455000 11.875000 2.465000 ;
        RECT 11.665000 0.825000 11.875000 1.455000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.200000 0.255000 10.485000 0.715000 ;
        RECT 10.200000 1.630000 10.485000 2.465000 ;
        RECT 10.305000 0.715000 10.485000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.235000 1.095000 9.690000 1.325000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.585000 0.735000 3.995000 0.965000 ;
        RECT 3.585000 0.965000 3.915000 1.065000 ;
      LAYER mcon ;
        RECT 3.825000 0.765000 3.995000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.280000 0.735000 7.825000 1.065000 ;
      LAYER mcon ;
        RECT 7.575000 0.765000 7.745000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765000 0.735000 4.055000 0.780000 ;
        RECT 3.765000 0.780000 7.805000 0.920000 ;
        RECT 3.765000 0.920000 4.055000 0.965000 ;
        RECT 7.515000 0.735000 7.805000 0.780000 ;
        RECT 7.515000 0.920000 7.805000 0.965000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.435000 1.625000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.150000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.840000 0.805000 ;
      RECT  0.175000  1.795000  0.840000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.610000  0.805000  0.840000 1.795000 ;
      RECT  1.015000  0.345000  1.235000 2.465000 ;
      RECT  1.405000  0.635000  2.125000 0.825000 ;
      RECT  1.405000  0.825000  1.575000 1.795000 ;
      RECT  1.405000  1.795000  2.125000 1.965000 ;
      RECT  1.430000  0.085000  1.785000 0.465000 ;
      RECT  1.430000  2.135000  1.785000 2.635000 ;
      RECT  1.955000  0.305000  2.125000 0.635000 ;
      RECT  1.955000  1.965000  2.125000 2.465000 ;
      RECT  2.325000  0.705000  2.545000 1.575000 ;
      RECT  2.325000  1.575000  2.825000 1.955000 ;
      RECT  2.335000  2.250000  3.165000 2.420000 ;
      RECT  2.400000  0.265000  3.415000 0.465000 ;
      RECT  2.725000  0.645000  3.075000 1.015000 ;
      RECT  2.995000  1.195000  3.415000 1.235000 ;
      RECT  2.995000  1.235000  4.345000 1.405000 ;
      RECT  2.995000  1.405000  3.165000 2.250000 ;
      RECT  3.245000  0.465000  3.415000 1.195000 ;
      RECT  3.335000  1.575000  3.585000 1.785000 ;
      RECT  3.335000  1.785000  4.685000 2.035000 ;
      RECT  3.405000  2.205000  3.785000 2.635000 ;
      RECT  3.585000  0.085000  3.755000 0.525000 ;
      RECT  3.925000  0.255000  5.075000 0.425000 ;
      RECT  3.925000  0.425000  4.255000 0.505000 ;
      RECT  4.085000  2.035000  4.255000 2.375000 ;
      RECT  4.095000  1.405000  4.345000 1.485000 ;
      RECT  4.125000  1.155000  4.345000 1.235000 ;
      RECT  4.405000  0.595000  4.735000 0.765000 ;
      RECT  4.515000  0.765000  4.735000 0.895000 ;
      RECT  4.515000  0.895000  5.825000 1.065000 ;
      RECT  4.515000  1.065000  4.685000 1.785000 ;
      RECT  4.855000  1.235000  5.185000 1.415000 ;
      RECT  4.855000  1.415000  5.860000 1.655000 ;
      RECT  4.875000  1.915000  5.205000 2.635000 ;
      RECT  4.905000  0.425000  5.075000 0.715000 ;
      RECT  5.325000  0.085000  5.675000 0.465000 ;
      RECT  5.495000  1.065000  5.825000 1.235000 ;
      RECT  6.060000  1.575000  6.295000 1.985000 ;
      RECT  6.065000  1.060000  6.405000 1.125000 ;
      RECT  6.065000  1.125000  6.740000 1.305000 ;
      RECT  6.185000  0.705000  6.405000 1.060000 ;
      RECT  6.250000  2.250000  7.080000 2.420000 ;
      RECT  6.300000  0.265000  7.080000 0.465000 ;
      RECT  6.535000  1.305000  6.740000 1.905000 ;
      RECT  6.910000  0.465000  7.080000 1.235000 ;
      RECT  6.910000  1.235000  8.260000 1.405000 ;
      RECT  6.910000  1.405000  7.080000 2.250000 ;
      RECT  7.250000  0.085000  7.575000 0.525000 ;
      RECT  7.250000  1.575000  7.500000 1.915000 ;
      RECT  7.250000  1.915000 10.030000 2.085000 ;
      RECT  7.320000  2.255000  7.700000 2.635000 ;
      RECT  7.745000  0.255000  8.955000 0.425000 ;
      RECT  7.745000  0.425000  8.075000 0.545000 ;
      RECT  7.940000  2.085000  8.110000 2.375000 ;
      RECT  8.040000  1.075000  8.260000 1.235000 ;
      RECT  8.215000  0.665000  8.615000 0.835000 ;
      RECT  8.430000  0.835000  8.615000 0.840000 ;
      RECT  8.430000  0.840000  8.600000 1.915000 ;
      RECT  8.640000  2.255000 10.030000 2.635000 ;
      RECT  8.770000  1.110000  9.055000 1.575000 ;
      RECT  8.770000  1.575000  9.555000 1.745000 ;
      RECT  8.785000  0.425000  8.955000 0.585000 ;
      RECT  8.835000  0.755000  9.475000 0.925000 ;
      RECT  8.835000  0.925000  9.055000 1.110000 ;
      RECT  9.265000  0.265000  9.475000 0.755000 ;
      RECT  9.725000  0.085000 10.030000 0.805000 ;
      RECT  9.860000  0.995000 10.125000 1.325000 ;
      RECT  9.860000  1.325000 10.030000 1.915000 ;
      RECT 10.660000  0.255000 10.975000 0.995000 ;
      RECT 10.660000  0.995000 11.495000 1.325000 ;
      RECT 10.660000  1.325000 10.975000 2.415000 ;
      RECT 11.150000  0.085000 11.445000 0.545000 ;
      RECT 11.155000  1.765000 11.445000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.610000  0.765000  0.780000 0.935000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  1.785000  1.235000 1.955000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  1.785000  2.615000 1.955000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  0.765000  3.075000 0.935000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  1.445000  5.835000 1.615000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  1.105000  6.295000 1.275000 ;
      RECT  6.125000  1.785000  6.295000 1.955000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.855000  1.445000  9.025000 1.615000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 0.735000 0.840000 0.780000 ;
      RECT 0.550000 0.780000 3.135000 0.920000 ;
      RECT 0.550000 0.920000 0.840000 0.965000 ;
      RECT 1.005000 1.755000 1.295000 1.800000 ;
      RECT 1.005000 1.800000 6.355000 1.940000 ;
      RECT 1.005000 1.940000 1.295000 1.985000 ;
      RECT 2.385000 1.755000 2.675000 1.800000 ;
      RECT 2.385000 1.940000 2.675000 1.985000 ;
      RECT 2.845000 0.735000 3.135000 0.780000 ;
      RECT 2.845000 0.920000 3.135000 0.965000 ;
      RECT 2.920000 0.965000 3.135000 1.120000 ;
      RECT 2.920000 1.120000 6.355000 1.260000 ;
      RECT 5.605000 1.415000 5.895000 1.460000 ;
      RECT 5.605000 1.460000 9.085000 1.600000 ;
      RECT 5.605000 1.600000 5.895000 1.645000 ;
      RECT 6.065000 1.075000 6.355000 1.120000 ;
      RECT 6.065000 1.260000 6.355000 1.305000 ;
      RECT 6.065000 1.755000 6.355000 1.800000 ;
      RECT 6.065000 1.940000 6.355000 1.985000 ;
      RECT 8.795000 1.415000 9.085000 1.460000 ;
      RECT 8.795000 1.600000 9.085000 1.645000 ;
  END
END sky130_fd_sc_hd__dfbbn_1
MACRO sky130_fd_sc_hd__dfbbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfbbn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.88000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.760000 1.005000 2.170000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.115000 0.255000 12.345000 0.825000 ;
        RECT 12.115000 1.445000 12.345000 2.465000 ;
        RECT 12.160000 0.825000 12.345000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.240000 0.255000 10.500000 0.715000 ;
        RECT 10.240000 1.630000 10.500000 2.465000 ;
        RECT 10.320000 0.715000 10.500000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.250000 1.095000 9.730000 1.325000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.600000 0.735000 4.010000 0.965000 ;
        RECT 3.600000 0.965000 3.930000 1.065000 ;
      LAYER mcon ;
        RECT 3.840000 0.765000 4.010000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.470000 0.735000 7.845000 1.065000 ;
      LAYER mcon ;
        RECT 7.520000 0.765000 7.690000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.780000 0.735000 4.070000 0.780000 ;
        RECT 3.780000 0.780000 7.750000 0.920000 ;
        RECT 3.780000 0.920000 4.070000 0.965000 ;
        RECT 7.460000 0.735000 7.750000 0.780000 ;
        RECT 7.460000 0.920000 7.750000 0.965000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.440000 1.625000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.880000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 13.070000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.880000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.880000 0.085000 ;
      RECT  0.000000  2.635000 12.880000 2.805000 ;
      RECT  0.085000  0.345000  0.345000 0.635000 ;
      RECT  0.085000  0.635000  0.840000 0.805000 ;
      RECT  0.085000  1.795000  0.840000 1.965000 ;
      RECT  0.085000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.610000  0.805000  0.840000 1.795000 ;
      RECT  1.015000  0.345000  1.240000 2.465000 ;
      RECT  1.420000  0.635000  2.125000 0.825000 ;
      RECT  1.420000  0.825000  1.590000 1.795000 ;
      RECT  1.420000  1.795000  2.125000 1.965000 ;
      RECT  1.445000  0.085000  1.785000 0.465000 ;
      RECT  1.445000  2.135000  1.785000 2.635000 ;
      RECT  1.955000  0.305000  2.125000 0.635000 ;
      RECT  1.955000  1.965000  2.125000 2.465000 ;
      RECT  2.340000  0.705000  2.560000 1.575000 ;
      RECT  2.340000  1.575000  2.840000 1.955000 ;
      RECT  2.350000  2.250000  3.180000 2.420000 ;
      RECT  2.415000  0.265000  3.410000 0.465000 ;
      RECT  2.740000  0.645000  3.070000 1.015000 ;
      RECT  3.010000  1.195000  3.410000 1.235000 ;
      RECT  3.010000  1.235000  4.360000 1.405000 ;
      RECT  3.010000  1.405000  3.180000 2.250000 ;
      RECT  3.240000  0.465000  3.410000 1.195000 ;
      RECT  3.350000  1.575000  3.600000 1.785000 ;
      RECT  3.350000  1.785000  4.700000 2.035000 ;
      RECT  3.420000  2.205000  3.800000 2.635000 ;
      RECT  3.580000  0.085000  3.750000 0.525000 ;
      RECT  3.920000  0.255000  5.170000 0.425000 ;
      RECT  3.920000  0.425000  4.250000 0.545000 ;
      RECT  4.100000  2.035000  4.270000 2.375000 ;
      RECT  4.110000  1.405000  4.360000 1.485000 ;
      RECT  4.140000  1.155000  4.360000 1.235000 ;
      RECT  4.420000  0.595000  4.750000 0.765000 ;
      RECT  4.530000  0.765000  4.750000 0.895000 ;
      RECT  4.530000  0.895000  5.840000 1.065000 ;
      RECT  4.530000  1.065000  4.700000 1.785000 ;
      RECT  4.870000  1.235000  5.200000 1.415000 ;
      RECT  4.870000  1.415000  5.875000 1.655000 ;
      RECT  4.890000  1.915000  5.220000 2.635000 ;
      RECT  4.920000  0.425000  5.170000 0.715000 ;
      RECT  5.360000  0.085000  5.690000 0.465000 ;
      RECT  5.510000  1.065000  5.840000 1.235000 ;
      RECT  6.075000  1.575000  6.310000 1.985000 ;
      RECT  6.135000  0.705000  6.420000 1.125000 ;
      RECT  6.135000  1.125000  6.755000 1.305000 ;
      RECT  6.265000  2.250000  7.095000 2.420000 ;
      RECT  6.330000  0.265000  7.095000 0.465000 ;
      RECT  6.550000  1.305000  6.755000 1.905000 ;
      RECT  6.925000  0.465000  7.095000 1.235000 ;
      RECT  6.925000  1.235000  8.275000 1.405000 ;
      RECT  6.925000  1.405000  7.095000 2.250000 ;
      RECT  7.265000  1.575000  7.515000 1.915000 ;
      RECT  7.265000  1.915000 10.070000 2.085000 ;
      RECT  7.275000  0.085000  7.535000 0.525000 ;
      RECT  7.335000  2.255000  7.715000 2.635000 ;
      RECT  7.795000  0.255000  8.965000 0.425000 ;
      RECT  7.795000  0.425000  8.125000 0.545000 ;
      RECT  7.955000  2.085000  8.125000 2.375000 ;
      RECT  8.055000  1.075000  8.275000 1.235000 ;
      RECT  8.295000  0.595000  8.625000 0.780000 ;
      RECT  8.445000  0.780000  8.625000 1.915000 ;
      RECT  8.655000  2.255000 10.070000 2.635000 ;
      RECT  8.795000  0.425000  8.965000 0.585000 ;
      RECT  8.795000  0.755000  9.500000 0.925000 ;
      RECT  8.795000  0.925000  9.070000 1.575000 ;
      RECT  8.795000  1.575000  9.570000 1.745000 ;
      RECT  9.280000  0.265000  9.500000 0.755000 ;
      RECT  9.740000  0.085000 10.070000 0.805000 ;
      RECT  9.900000  0.995000 10.140000 1.325000 ;
      RECT  9.900000  1.325000 10.070000 1.915000 ;
      RECT 10.680000  0.085000 10.910000 0.885000 ;
      RECT 10.680000  1.465000 10.910000 2.635000 ;
      RECT 11.215000  0.255000 11.470000 0.995000 ;
      RECT 11.215000  0.995000 11.990000 1.325000 ;
      RECT 11.215000  1.325000 11.470000 2.415000 ;
      RECT 11.650000  0.085000 11.945000 0.545000 ;
      RECT 11.650000  1.765000 11.945000 2.635000 ;
      RECT 12.515000  0.085000 12.795000 0.885000 ;
      RECT 12.515000  1.465000 12.795000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.610000  0.765000  0.780000 0.935000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.070000  1.785000  1.240000 1.955000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.460000  1.785000  2.630000 1.955000 ;
      RECT  2.900000  0.765000  3.070000 0.935000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.680000  1.445000  5.850000 1.615000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.140000  1.105000  6.310000 1.275000 ;
      RECT  6.140000  1.785000  6.310000 1.955000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  8.900000  1.445000  9.070000 1.615000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 0.735000 0.840000 0.780000 ;
      RECT 0.550000 0.780000 3.130000 0.920000 ;
      RECT 0.550000 0.920000 0.840000 0.965000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 6.370000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.400000 1.755000 2.690000 1.800000 ;
      RECT 2.400000 1.940000 2.690000 1.985000 ;
      RECT 2.840000 0.735000 3.130000 0.780000 ;
      RECT 2.840000 0.920000 3.130000 0.965000 ;
      RECT 2.935000 0.965000 3.130000 1.120000 ;
      RECT 2.935000 1.120000 6.370000 1.260000 ;
      RECT 5.620000 1.415000 5.910000 1.460000 ;
      RECT 5.620000 1.460000 9.130000 1.600000 ;
      RECT 5.620000 1.600000 5.910000 1.645000 ;
      RECT 6.080000 1.075000 6.370000 1.120000 ;
      RECT 6.080000 1.260000 6.370000 1.305000 ;
      RECT 6.080000 1.755000 6.370000 1.800000 ;
      RECT 6.080000 1.940000 6.370000 1.985000 ;
      RECT 8.840000 1.415000 9.130000 1.460000 ;
      RECT 8.840000 1.600000 9.130000 1.645000 ;
  END
END sky130_fd_sc_hd__dfbbn_2
MACRO sky130_fd_sc_hd__dfbbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfbbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.750000 1.005000 2.160000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.615000 0.255000 11.875000 0.825000 ;
        RECT 11.615000 1.445000 11.875000 2.465000 ;
        RECT 11.660000 0.825000 11.875000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.200000 0.255000 10.485000 0.715000 ;
        RECT 10.200000 1.630000 10.485000 2.465000 ;
        RECT 10.280000 0.715000 10.485000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.315000 1.095000 9.690000 1.325000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.590000 0.735000 4.000000 0.965000 ;
        RECT 3.590000 0.965000 3.920000 1.065000 ;
      LAYER mcon ;
        RECT 3.830000 0.765000 4.000000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.460000 0.735000 7.835000 1.065000 ;
      LAYER mcon ;
        RECT 7.510000 0.765000 7.680000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.770000 0.735000 4.060000 0.780000 ;
        RECT 3.770000 0.780000 7.740000 0.920000 ;
        RECT 3.770000 0.920000 4.060000 0.965000 ;
        RECT 7.450000 0.735000 7.740000 0.780000 ;
        RECT 7.450000 0.920000 7.740000 0.965000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.150000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.085000  0.345000  0.345000 0.635000 ;
      RECT  0.085000  0.635000  0.840000 0.805000 ;
      RECT  0.085000  1.795000  0.840000 1.965000 ;
      RECT  0.085000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.610000  0.805000  0.840000 1.795000 ;
      RECT  1.015000  0.345000  1.240000 2.465000 ;
      RECT  1.410000  0.635000  2.125000 0.825000 ;
      RECT  1.410000  0.825000  1.580000 1.795000 ;
      RECT  1.410000  1.795000  2.125000 1.965000 ;
      RECT  1.435000  0.085000  1.785000 0.465000 ;
      RECT  1.435000  2.135000  1.785000 2.635000 ;
      RECT  1.955000  0.305000  2.125000 0.635000 ;
      RECT  1.955000  1.965000  2.125000 2.465000 ;
      RECT  2.330000  0.705000  2.550000 1.575000 ;
      RECT  2.330000  1.575000  2.830000 1.955000 ;
      RECT  2.340000  2.250000  3.170000 2.420000 ;
      RECT  2.405000  0.265000  3.400000 0.465000 ;
      RECT  2.730000  0.645000  3.060000 1.015000 ;
      RECT  3.000000  1.195000  3.400000 1.235000 ;
      RECT  3.000000  1.235000  4.350000 1.405000 ;
      RECT  3.000000  1.405000  3.170000 2.250000 ;
      RECT  3.230000  0.465000  3.400000 1.195000 ;
      RECT  3.340000  1.575000  3.590000 1.785000 ;
      RECT  3.340000  1.785000  4.690000 2.035000 ;
      RECT  3.410000  2.205000  3.790000 2.635000 ;
      RECT  3.570000  0.085000  3.740000 0.525000 ;
      RECT  3.910000  0.255000  5.080000 0.425000 ;
      RECT  3.910000  0.425000  4.240000 0.545000 ;
      RECT  4.090000  2.035000  4.260000 2.375000 ;
      RECT  4.100000  1.405000  4.350000 1.485000 ;
      RECT  4.130000  1.155000  4.350000 1.235000 ;
      RECT  4.410000  0.595000  4.740000 0.765000 ;
      RECT  4.520000  0.765000  4.740000 0.895000 ;
      RECT  4.520000  0.895000  5.830000 1.065000 ;
      RECT  4.520000  1.065000  4.690000 1.785000 ;
      RECT  4.860000  1.235000  5.190000 1.415000 ;
      RECT  4.860000  1.415000  5.865000 1.655000 ;
      RECT  4.880000  1.915000  5.210000 2.635000 ;
      RECT  4.910000  0.425000  5.080000 0.715000 ;
      RECT  5.350000  0.085000  5.680000 0.465000 ;
      RECT  5.500000  1.065000  5.830000 1.235000 ;
      RECT  6.065000  1.575000  6.300000 1.985000 ;
      RECT  6.125000  0.705000  6.410000 1.125000 ;
      RECT  6.125000  1.125000  6.745000 1.305000 ;
      RECT  6.255000  2.250000  7.085000 2.420000 ;
      RECT  6.320000  0.265000  7.085000 0.465000 ;
      RECT  6.540000  1.305000  6.745000 1.905000 ;
      RECT  6.915000  0.465000  7.085000 1.235000 ;
      RECT  6.915000  1.235000  8.265000 1.405000 ;
      RECT  6.915000  1.405000  7.085000 2.250000 ;
      RECT  7.255000  1.575000  7.505000 1.915000 ;
      RECT  7.255000  1.915000 10.030000 2.085000 ;
      RECT  7.265000  0.085000  7.525000 0.525000 ;
      RECT  7.325000  2.255000  7.705000 2.635000 ;
      RECT  7.785000  0.255000  8.955000 0.425000 ;
      RECT  7.785000  0.425000  8.115000 0.545000 ;
      RECT  7.945000  2.085000  8.115000 2.375000 ;
      RECT  8.045000  1.075000  8.265000 1.235000 ;
      RECT  8.285000  0.595000  8.615000 0.780000 ;
      RECT  8.435000  0.780000  8.615000 1.915000 ;
      RECT  8.645000  2.255000 10.030000 2.635000 ;
      RECT  8.785000  0.425000  8.955000 0.585000 ;
      RECT  8.785000  0.755000  9.475000 0.925000 ;
      RECT  8.785000  0.925000  9.060000 1.575000 ;
      RECT  8.785000  1.575000  9.545000 1.745000 ;
      RECT  9.240000  0.265000  9.475000 0.755000 ;
      RECT  9.700000  0.085000 10.030000 0.805000 ;
      RECT  9.860000  0.995000 10.110000 1.325000 ;
      RECT  9.860000  1.325000 10.030000 1.915000 ;
      RECT 10.655000  0.255000 10.970000 0.995000 ;
      RECT 10.655000  0.995000 11.490000 1.325000 ;
      RECT 10.655000  1.325000 10.970000 2.415000 ;
      RECT 11.150000  0.085000 11.445000 0.545000 ;
      RECT 11.150000  1.765000 11.445000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.610000  1.785000  0.780000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.070000  0.765000  1.240000 0.935000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.450000  1.785000  2.620000 1.955000 ;
      RECT  2.890000  0.765000  3.060000 0.935000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.670000  1.445000  5.840000 1.615000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.130000  1.105000  6.300000 1.275000 ;
      RECT  6.130000  1.785000  6.300000 1.955000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  8.890000  1.445000  9.060000 1.615000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.755000 0.840000 1.800000 ;
      RECT 0.550000 1.800000 6.360000 1.940000 ;
      RECT 0.550000 1.940000 0.840000 1.985000 ;
      RECT 1.010000 0.735000 1.300000 0.780000 ;
      RECT 1.010000 0.780000 3.120000 0.920000 ;
      RECT 1.010000 0.920000 1.300000 0.965000 ;
      RECT 2.390000 1.755000 2.680000 1.800000 ;
      RECT 2.390000 1.940000 2.680000 1.985000 ;
      RECT 2.830000 0.735000 3.120000 0.780000 ;
      RECT 2.830000 0.920000 3.120000 0.965000 ;
      RECT 2.925000 0.965000 3.120000 1.120000 ;
      RECT 2.925000 1.120000 6.360000 1.260000 ;
      RECT 5.610000 1.415000 5.900000 1.460000 ;
      RECT 5.610000 1.460000 9.120000 1.600000 ;
      RECT 5.610000 1.600000 5.900000 1.645000 ;
      RECT 6.070000 1.075000 6.360000 1.120000 ;
      RECT 6.070000 1.260000 6.360000 1.305000 ;
      RECT 6.070000 1.755000 6.360000 1.800000 ;
      RECT 6.070000 1.940000 6.360000 1.985000 ;
      RECT 8.830000 1.415000 9.120000 1.460000 ;
      RECT 8.830000 1.600000 9.120000 1.645000 ;
  END
END sky130_fd_sc_hd__dfbbp_1
MACRO sky130_fd_sc_hd__dfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.58000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.665000 1.680000 2.450000 ;
        RECT 1.415000 0.615000 1.875000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.600000 1.455000 9.005000 2.465000 ;
        RECT 8.675000 0.275000 9.005000 1.455000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.180000 0.265000 10.435000 0.795000 ;
        RECT 10.180000 1.445000 10.435000 2.325000 ;
        RECT 10.225000 0.795000 10.435000 1.445000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.765000 4.595000 1.015000 ;
      LAYER mcon ;
        RECT 4.165000 0.765000 4.335000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105000 1.035000 7.645000 1.405000 ;
        RECT 7.405000 0.635000 7.645000 1.035000 ;
      LAYER mcon ;
        RECT 7.105000 1.080000 7.275000 1.250000 ;
        RECT 7.405000 0.765000 7.575000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745000 0.735000 4.395000 0.780000 ;
        RECT 3.745000 0.780000 7.635000 0.920000 ;
        RECT 3.745000 0.920000 4.395000 0.965000 ;
        RECT 7.045000 0.920000 7.635000 0.965000 ;
        RECT 7.045000 0.965000 7.335000 1.280000 ;
        RECT 7.345000 0.735000 7.635000 0.780000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.770000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.580000 0.085000 ;
      RECT 0.000000  2.635000 10.580000 2.805000 ;
      RECT 0.090000  0.345000  0.345000 0.635000 ;
      RECT 0.090000  0.635000  0.840000 0.805000 ;
      RECT 0.090000  1.795000  0.840000 1.965000 ;
      RECT 0.090000  1.965000  0.345000 2.465000 ;
      RECT 0.515000  0.085000  0.845000 0.465000 ;
      RECT 0.515000  2.135000  0.845000 2.635000 ;
      RECT 0.610000  0.805000  0.840000 1.795000 ;
      RECT 1.015000  0.345000  1.185000 2.465000 ;
      RECT 1.545000  0.085000  1.875000 0.445000 ;
      RECT 1.850000  2.175000  2.100000 2.635000 ;
      RECT 2.045000  0.305000  2.540000 0.475000 ;
      RECT 2.045000  0.475000  2.215000 1.835000 ;
      RECT 2.045000  1.835000  2.440000 2.005000 ;
      RECT 2.270000  2.005000  2.440000 2.135000 ;
      RECT 2.270000  2.135000  2.520000 2.465000 ;
      RECT 2.385000  0.765000  2.735000 1.385000 ;
      RECT 2.610000  1.575000  3.075000 1.965000 ;
      RECT 2.735000  2.135000  3.415000 2.465000 ;
      RECT 2.745000  0.305000  3.600000 0.475000 ;
      RECT 2.905000  0.765000  3.260000 0.985000 ;
      RECT 2.905000  0.985000  3.075000 1.575000 ;
      RECT 3.245000  1.185000  4.935000 1.355000 ;
      RECT 3.245000  1.355000  3.415000 2.135000 ;
      RECT 3.430000  0.475000  3.600000 1.185000 ;
      RECT 3.585000  1.865000  4.660000 2.035000 ;
      RECT 3.585000  2.035000  3.755000 2.375000 ;
      RECT 3.775000  1.525000  5.275000 1.695000 ;
      RECT 3.990000  2.205000  4.320000 2.635000 ;
      RECT 4.475000  0.085000  4.805000 0.545000 ;
      RECT 4.490000  2.035000  4.660000 2.375000 ;
      RECT 4.765000  1.005000  4.935000 1.185000 ;
      RECT 4.955000  2.175000  5.325000 2.635000 ;
      RECT 5.015000  0.275000  5.365000 0.445000 ;
      RECT 5.015000  0.445000  5.275000 0.835000 ;
      RECT 5.105000  0.835000  5.275000 1.525000 ;
      RECT 5.105000  1.695000  5.275000 1.835000 ;
      RECT 5.105000  1.835000  5.665000 2.005000 ;
      RECT 5.465000  0.705000  5.675000 1.495000 ;
      RECT 5.465000  1.495000  6.140000 1.655000 ;
      RECT 5.465000  1.655000  6.430000 1.665000 ;
      RECT 5.495000  2.005000  5.665000 2.465000 ;
      RECT 5.585000  0.255000  6.535000 0.535000 ;
      RECT 5.845000  0.705000  6.195000 1.325000 ;
      RECT 5.900000  2.125000  6.770000 2.465000 ;
      RECT 5.970000  1.665000  6.430000 1.955000 ;
      RECT 6.365000  0.535000  6.535000 1.315000 ;
      RECT 6.365000  1.315000  6.770000 1.485000 ;
      RECT 6.600000  1.485000  6.770000 1.575000 ;
      RECT 6.600000  1.575000  7.820000 1.745000 ;
      RECT 6.600000  1.745000  6.770000 2.125000 ;
      RECT 6.705000  0.085000  6.895000 0.525000 ;
      RECT 6.705000  0.695000  7.235000 0.865000 ;
      RECT 6.705000  0.865000  6.925000 1.145000 ;
      RECT 6.940000  2.175000  7.190000 2.635000 ;
      RECT 7.065000  0.295000  8.135000 0.465000 ;
      RECT 7.065000  0.465000  7.235000 0.695000 ;
      RECT 7.360000  1.915000  8.160000 2.085000 ;
      RECT 7.360000  2.085000  7.530000 2.375000 ;
      RECT 7.710000  2.255000  8.430000 2.635000 ;
      RECT 7.815000  0.465000  8.135000 0.820000 ;
      RECT 7.815000  0.820000  8.140000 0.995000 ;
      RECT 7.815000  0.995000  8.435000 1.295000 ;
      RECT 7.990000  1.295000  8.435000 1.325000 ;
      RECT 7.990000  1.325000  8.160000 1.915000 ;
      RECT 8.335000  0.085000  8.505000 0.770000 ;
      RECT 9.195000  0.345000  9.445000 0.995000 ;
      RECT 9.195000  0.995000 10.055000 1.325000 ;
      RECT 9.195000  1.325000  9.525000 2.425000 ;
      RECT 9.760000  0.085000  9.930000 0.680000 ;
      RECT 9.760000  1.495000  9.930000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.610000  1.105000  0.780000 1.275000 ;
      RECT  1.015000  1.785000  1.185000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  1.105000  2.615000 1.275000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  1.785000  3.075000 1.955000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.025000  1.105000  6.195000 1.275000 ;
      RECT  6.025000  1.785000  6.195000 1.955000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.075000 0.840000 1.120000 ;
      RECT 0.550000 1.120000 6.255000 1.260000 ;
      RECT 0.550000 1.260000 0.840000 1.305000 ;
      RECT 0.955000 1.755000 1.245000 1.800000 ;
      RECT 0.955000 1.800000 6.255000 1.940000 ;
      RECT 0.955000 1.940000 1.245000 1.985000 ;
      RECT 2.385000 1.075000 2.675000 1.120000 ;
      RECT 2.385000 1.260000 2.675000 1.305000 ;
      RECT 2.845000 1.755000 3.135000 1.800000 ;
      RECT 2.845000 1.940000 3.135000 1.985000 ;
      RECT 5.965000 1.075000 6.255000 1.120000 ;
      RECT 5.965000 1.260000 6.255000 1.305000 ;
      RECT 5.965000 1.755000 6.255000 1.800000 ;
      RECT 5.965000 1.940000 6.255000 1.985000 ;
  END
END sky130_fd_sc_hd__dfrbp_1
MACRO sky130_fd_sc_hd__dfrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.665000 1.680000 2.450000 ;
        RECT 1.415000 0.615000 1.875000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.160000 0.265000 9.495000 1.695000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.030000 1.535000 10.420000 2.080000 ;
        RECT 10.040000 0.310000 10.420000 0.825000 ;
        RECT 10.120000 2.080000 10.420000 2.465000 ;
        RECT 10.250000 0.825000 10.420000 1.535000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.765000 4.595000 1.015000 ;
      LAYER mcon ;
        RECT 4.165000 0.765000 4.335000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105000 1.035000 7.645000 1.405000 ;
        RECT 7.405000 0.635000 7.645000 1.035000 ;
      LAYER mcon ;
        RECT 7.105000 1.080000 7.275000 1.250000 ;
        RECT 7.405000 0.765000 7.575000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745000 0.735000 4.395000 0.780000 ;
        RECT 3.745000 0.780000 7.635000 0.920000 ;
        RECT 3.745000 0.920000 4.395000 0.965000 ;
        RECT 7.045000 0.920000 7.635000 0.965000 ;
        RECT 7.045000 0.965000 7.335000 1.280000 ;
        RECT 7.345000 0.735000 7.635000 0.780000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.090000  0.345000  0.345000 0.635000 ;
      RECT  0.090000  0.635000  0.840000 0.805000 ;
      RECT  0.090000  1.795000  0.840000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.610000  0.805000  0.840000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.545000  0.085000  1.875000 0.445000 ;
      RECT  1.850000  2.175000  2.100000 2.635000 ;
      RECT  2.045000  0.305000  2.540000 0.475000 ;
      RECT  2.045000  0.475000  2.215000 1.835000 ;
      RECT  2.045000  1.835000  2.440000 2.005000 ;
      RECT  2.270000  2.005000  2.440000 2.135000 ;
      RECT  2.270000  2.135000  2.520000 2.465000 ;
      RECT  2.385000  0.765000  2.735000 1.385000 ;
      RECT  2.610000  1.575000  3.075000 1.965000 ;
      RECT  2.735000  2.135000  3.415000 2.465000 ;
      RECT  2.745000  0.305000  3.600000 0.475000 ;
      RECT  2.905000  0.765000  3.260000 0.985000 ;
      RECT  2.905000  0.985000  3.075000 1.575000 ;
      RECT  3.245000  1.185000  4.935000 1.355000 ;
      RECT  3.245000  1.355000  3.415000 2.135000 ;
      RECT  3.430000  0.475000  3.600000 1.185000 ;
      RECT  3.585000  1.865000  4.660000 2.035000 ;
      RECT  3.585000  2.035000  3.755000 2.375000 ;
      RECT  3.775000  1.525000  5.275000 1.695000 ;
      RECT  3.990000  2.205000  4.320000 2.635000 ;
      RECT  4.475000  0.085000  4.805000 0.545000 ;
      RECT  4.490000  2.035000  4.660000 2.375000 ;
      RECT  4.765000  1.005000  4.935000 1.185000 ;
      RECT  4.955000  2.175000  5.325000 2.635000 ;
      RECT  5.015000  0.275000  5.365000 0.445000 ;
      RECT  5.015000  0.445000  5.275000 0.835000 ;
      RECT  5.105000  0.835000  5.275000 1.525000 ;
      RECT  5.105000  1.695000  5.275000 1.835000 ;
      RECT  5.105000  1.835000  5.665000 2.005000 ;
      RECT  5.465000  0.705000  5.675000 1.495000 ;
      RECT  5.465000  1.495000  6.140000 1.655000 ;
      RECT  5.465000  1.655000  6.430000 1.665000 ;
      RECT  5.495000  2.005000  5.665000 2.465000 ;
      RECT  5.585000  0.255000  6.535000 0.535000 ;
      RECT  5.845000  0.705000  6.195000 1.325000 ;
      RECT  5.900000  2.125000  6.770000 2.465000 ;
      RECT  5.970000  1.665000  6.430000 1.955000 ;
      RECT  6.365000  0.535000  6.535000 1.315000 ;
      RECT  6.365000  1.315000  6.770000 1.485000 ;
      RECT  6.600000  1.485000  6.770000 1.575000 ;
      RECT  6.600000  1.575000  7.820000 1.745000 ;
      RECT  6.600000  1.745000  6.770000 2.125000 ;
      RECT  6.705000  0.085000  6.895000 0.525000 ;
      RECT  6.705000  0.695000  7.235000 0.865000 ;
      RECT  6.705000  0.865000  6.925000 1.145000 ;
      RECT  6.940000  2.175000  7.190000 2.635000 ;
      RECT  7.065000  0.295000  7.985000 0.465000 ;
      RECT  7.065000  0.465000  7.235000 0.695000 ;
      RECT  7.360000  1.915000  8.160000 2.085000 ;
      RECT  7.360000  2.085000  7.530000 2.375000 ;
      RECT  7.710000  2.255000  8.055000 2.635000 ;
      RECT  7.815000  0.465000  7.985000 0.995000 ;
      RECT  7.815000  0.995000  8.160000 1.075000 ;
      RECT  7.815000  1.075000  8.650000 1.295000 ;
      RECT  7.990000  1.295000  8.650000 1.325000 ;
      RECT  7.990000  1.325000  8.160000 1.915000 ;
      RECT  8.335000  0.345000  8.585000 0.715000 ;
      RECT  8.335000  0.715000  8.990000 0.885000 ;
      RECT  8.335000  1.795000  8.990000 1.865000 ;
      RECT  8.335000  1.865000  9.835000 2.035000 ;
      RECT  8.335000  2.035000  8.560000 2.465000 ;
      RECT  8.730000  2.205000  9.070000 2.635000 ;
      RECT  8.755000  0.085000  8.990000 0.545000 ;
      RECT  8.820000  0.885000  8.990000 1.795000 ;
      RECT  9.620000  2.255000  9.950000 2.635000 ;
      RECT  9.665000  0.995000 10.080000 1.325000 ;
      RECT  9.665000  1.325000  9.835000 1.865000 ;
      RECT  9.700000  0.085000  9.870000 0.825000 ;
      RECT 10.590000  0.085000 10.760000 0.930000 ;
      RECT 10.590000  1.445000 10.760000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.610000  1.105000  0.780000 1.275000 ;
      RECT  1.015000  1.785000  1.185000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  1.105000  2.615000 1.275000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  1.785000  3.075000 1.955000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.025000  1.105000  6.195000 1.275000 ;
      RECT  6.025000  1.785000  6.195000 1.955000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.075000 0.840000 1.120000 ;
      RECT 0.550000 1.120000 6.255000 1.260000 ;
      RECT 0.550000 1.260000 0.840000 1.305000 ;
      RECT 0.955000 1.755000 1.245000 1.800000 ;
      RECT 0.955000 1.800000 6.255000 1.940000 ;
      RECT 0.955000 1.940000 1.245000 1.985000 ;
      RECT 2.385000 1.075000 2.675000 1.120000 ;
      RECT 2.385000 1.260000 2.675000 1.305000 ;
      RECT 2.845000 1.755000 3.135000 1.800000 ;
      RECT 2.845000 1.940000 3.135000 1.985000 ;
      RECT 5.965000 1.075000 6.255000 1.120000 ;
      RECT 5.965000 1.260000 6.255000 1.305000 ;
      RECT 5.965000 1.755000 6.255000 1.800000 ;
      RECT 5.965000 1.940000 6.255000 1.985000 ;
  END
END sky130_fd_sc_hd__dfrbp_2
MACRO sky130_fd_sc_hd__dfrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.665000 1.680000 2.450000 ;
        RECT 1.415000 0.615000 1.875000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.855000 0.265000 9.110000 0.795000 ;
        RECT 8.855000 1.445000 9.110000 2.325000 ;
        RECT 8.900000 0.795000 9.110000 1.445000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.765000 4.595000 1.015000 ;
      LAYER mcon ;
        RECT 4.165000 0.765000 4.335000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105000 1.035000 7.645000 1.405000 ;
        RECT 7.405000 0.635000 7.645000 1.035000 ;
      LAYER mcon ;
        RECT 7.105000 1.080000 7.275000 1.250000 ;
        RECT 7.405000 0.765000 7.575000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745000 0.735000 4.395000 0.780000 ;
        RECT 3.745000 0.780000 7.635000 0.920000 ;
        RECT 3.745000 0.920000 4.395000 0.965000 ;
        RECT 7.045000 0.920000 7.635000 0.965000 ;
        RECT 7.045000 0.965000 7.335000 1.280000 ;
        RECT 7.345000 0.735000 7.635000 0.780000 ;
    END
  END RESET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.090000  0.345000 0.345000 0.635000 ;
      RECT 0.090000  0.635000 0.840000 0.805000 ;
      RECT 0.090000  1.795000 0.840000 1.965000 ;
      RECT 0.090000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 2.465000 ;
      RECT 1.545000  0.085000 1.875000 0.445000 ;
      RECT 1.850000  2.175000 2.100000 2.635000 ;
      RECT 2.045000  0.305000 2.540000 0.475000 ;
      RECT 2.045000  0.475000 2.215000 1.835000 ;
      RECT 2.045000  1.835000 2.440000 2.005000 ;
      RECT 2.270000  2.005000 2.440000 2.135000 ;
      RECT 2.270000  2.135000 2.520000 2.465000 ;
      RECT 2.385000  0.765000 2.735000 1.385000 ;
      RECT 2.610000  1.575000 3.075000 1.965000 ;
      RECT 2.735000  2.135000 3.415000 2.465000 ;
      RECT 2.745000  0.305000 3.600000 0.475000 ;
      RECT 2.905000  0.765000 3.260000 0.985000 ;
      RECT 2.905000  0.985000 3.075000 1.575000 ;
      RECT 3.245000  1.185000 4.935000 1.355000 ;
      RECT 3.245000  1.355000 3.415000 2.135000 ;
      RECT 3.430000  0.475000 3.600000 1.185000 ;
      RECT 3.585000  1.865000 4.660000 2.035000 ;
      RECT 3.585000  2.035000 3.755000 2.375000 ;
      RECT 3.775000  1.525000 5.275000 1.695000 ;
      RECT 3.990000  2.205000 4.320000 2.635000 ;
      RECT 4.475000  0.085000 4.805000 0.545000 ;
      RECT 4.490000  2.035000 4.660000 2.375000 ;
      RECT 4.765000  1.005000 4.935000 1.185000 ;
      RECT 4.955000  2.175000 5.325000 2.635000 ;
      RECT 5.015000  0.275000 5.365000 0.445000 ;
      RECT 5.015000  0.445000 5.275000 0.835000 ;
      RECT 5.105000  0.835000 5.275000 1.525000 ;
      RECT 5.105000  1.695000 5.275000 1.835000 ;
      RECT 5.105000  1.835000 5.665000 2.005000 ;
      RECT 5.465000  0.705000 5.675000 1.495000 ;
      RECT 5.465000  1.495000 6.140000 1.655000 ;
      RECT 5.465000  1.655000 6.430000 1.665000 ;
      RECT 5.495000  2.005000 5.665000 2.465000 ;
      RECT 5.585000  0.255000 6.535000 0.535000 ;
      RECT 5.845000  0.705000 6.195000 1.325000 ;
      RECT 5.900000  2.125000 6.770000 2.465000 ;
      RECT 5.970000  1.665000 6.430000 1.955000 ;
      RECT 6.365000  0.535000 6.535000 1.315000 ;
      RECT 6.365000  1.315000 6.770000 1.485000 ;
      RECT 6.600000  1.485000 6.770000 1.575000 ;
      RECT 6.600000  1.575000 7.820000 1.745000 ;
      RECT 6.600000  1.745000 6.770000 2.125000 ;
      RECT 6.705000  0.085000 6.895000 0.525000 ;
      RECT 6.705000  0.695000 7.235000 0.865000 ;
      RECT 6.705000  0.865000 6.925000 1.145000 ;
      RECT 6.940000  2.175000 7.190000 2.635000 ;
      RECT 7.065000  0.295000 8.135000 0.465000 ;
      RECT 7.065000  0.465000 7.235000 0.695000 ;
      RECT 7.360000  1.915000 8.160000 2.085000 ;
      RECT 7.360000  2.085000 7.530000 2.375000 ;
      RECT 7.710000  2.255000 8.040000 2.635000 ;
      RECT 7.815000  0.465000 8.135000 0.820000 ;
      RECT 7.815000  0.820000 8.140000 0.995000 ;
      RECT 7.815000  0.995000 8.730000 1.295000 ;
      RECT 7.990000  1.295000 8.730000 1.325000 ;
      RECT 7.990000  1.325000 8.160000 1.915000 ;
      RECT 8.380000  0.085000 8.685000 0.545000 ;
      RECT 8.380000  1.495000 8.685000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.655000  1.785000 0.825000 1.955000 ;
      RECT 1.015000  1.105000 1.185000 1.275000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  1.105000 2.615000 1.275000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  1.785000 3.075000 1.955000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.025000  1.105000 6.195000 1.275000 ;
      RECT 6.025000  1.785000 6.195000 1.955000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
    LAYER met1 ;
      RECT 0.595000 1.755000 0.885000 1.800000 ;
      RECT 0.595000 1.800000 6.255000 1.940000 ;
      RECT 0.595000 1.940000 0.885000 1.985000 ;
      RECT 0.955000 1.075000 1.245000 1.120000 ;
      RECT 0.955000 1.120000 6.255000 1.260000 ;
      RECT 0.955000 1.260000 1.245000 1.305000 ;
      RECT 2.385000 1.075000 2.675000 1.120000 ;
      RECT 2.385000 1.260000 2.675000 1.305000 ;
      RECT 2.845000 1.755000 3.135000 1.800000 ;
      RECT 2.845000 1.940000 3.135000 1.985000 ;
      RECT 5.965000 1.075000 6.255000 1.120000 ;
      RECT 5.965000 1.260000 6.255000 1.305000 ;
      RECT 5.965000 1.755000 6.255000 1.800000 ;
      RECT 5.965000 1.940000 6.255000 1.985000 ;
  END
END sky130_fd_sc_hd__dfrtn_1
MACRO sky130_fd_sc_hd__dfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.665000 1.680000 2.450000 ;
        RECT 1.415000 0.615000 1.875000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.855000 0.265000 9.110000 0.795000 ;
        RECT 8.855000 1.445000 9.110000 2.325000 ;
        RECT 8.900000 0.795000 9.110000 1.445000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.765000 4.595000 1.015000 ;
      LAYER mcon ;
        RECT 4.165000 0.765000 4.335000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105000 1.035000 7.645000 1.405000 ;
        RECT 7.405000 0.635000 7.645000 1.035000 ;
      LAYER mcon ;
        RECT 7.105000 1.080000 7.275000 1.250000 ;
        RECT 7.405000 0.765000 7.575000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745000 0.735000 4.395000 0.780000 ;
        RECT 3.745000 0.780000 7.635000 0.920000 ;
        RECT 3.745000 0.920000 4.395000 0.965000 ;
        RECT 7.045000 0.920000 7.635000 0.965000 ;
        RECT 7.045000 0.965000 7.335000 1.280000 ;
        RECT 7.345000 0.735000 7.635000 0.780000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.090000  0.345000 0.345000 0.635000 ;
      RECT 0.090000  0.635000 0.840000 0.805000 ;
      RECT 0.090000  1.795000 0.840000 1.965000 ;
      RECT 0.090000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 2.465000 ;
      RECT 1.545000  0.085000 1.875000 0.445000 ;
      RECT 1.850000  2.175000 2.100000 2.635000 ;
      RECT 2.045000  0.305000 2.540000 0.475000 ;
      RECT 2.045000  0.475000 2.215000 1.835000 ;
      RECT 2.045000  1.835000 2.440000 2.005000 ;
      RECT 2.270000  2.005000 2.440000 2.135000 ;
      RECT 2.270000  2.135000 2.520000 2.465000 ;
      RECT 2.385000  0.765000 2.735000 1.385000 ;
      RECT 2.610000  1.575000 3.075000 1.965000 ;
      RECT 2.735000  2.135000 3.415000 2.465000 ;
      RECT 2.745000  0.305000 3.600000 0.475000 ;
      RECT 2.905000  0.765000 3.260000 0.985000 ;
      RECT 2.905000  0.985000 3.075000 1.575000 ;
      RECT 3.245000  1.185000 4.935000 1.355000 ;
      RECT 3.245000  1.355000 3.415000 2.135000 ;
      RECT 3.430000  0.475000 3.600000 1.185000 ;
      RECT 3.585000  1.865000 4.660000 2.035000 ;
      RECT 3.585000  2.035000 3.755000 2.375000 ;
      RECT 3.775000  1.525000 5.275000 1.695000 ;
      RECT 3.990000  2.205000 4.320000 2.635000 ;
      RECT 4.475000  0.085000 4.805000 0.545000 ;
      RECT 4.490000  2.035000 4.660000 2.375000 ;
      RECT 4.765000  1.005000 4.935000 1.185000 ;
      RECT 4.955000  2.175000 5.325000 2.635000 ;
      RECT 5.015000  0.275000 5.365000 0.445000 ;
      RECT 5.015000  0.445000 5.275000 0.835000 ;
      RECT 5.105000  0.835000 5.275000 1.525000 ;
      RECT 5.105000  1.695000 5.275000 1.835000 ;
      RECT 5.105000  1.835000 5.665000 2.005000 ;
      RECT 5.465000  0.705000 5.675000 1.495000 ;
      RECT 5.465000  1.495000 6.140000 1.655000 ;
      RECT 5.465000  1.655000 6.430000 1.665000 ;
      RECT 5.495000  2.005000 5.665000 2.465000 ;
      RECT 5.585000  0.255000 6.535000 0.535000 ;
      RECT 5.845000  0.705000 6.195000 1.325000 ;
      RECT 5.900000  2.125000 6.770000 2.465000 ;
      RECT 5.970000  1.665000 6.430000 1.955000 ;
      RECT 6.365000  0.535000 6.535000 1.315000 ;
      RECT 6.365000  1.315000 6.770000 1.485000 ;
      RECT 6.600000  1.485000 6.770000 1.575000 ;
      RECT 6.600000  1.575000 7.820000 1.745000 ;
      RECT 6.600000  1.745000 6.770000 2.125000 ;
      RECT 6.705000  0.085000 6.895000 0.525000 ;
      RECT 6.705000  0.695000 7.235000 0.865000 ;
      RECT 6.705000  0.865000 6.925000 1.145000 ;
      RECT 6.940000  2.175000 7.190000 2.635000 ;
      RECT 7.065000  0.295000 8.135000 0.465000 ;
      RECT 7.065000  0.465000 7.235000 0.695000 ;
      RECT 7.360000  1.915000 8.160000 2.085000 ;
      RECT 7.360000  2.085000 7.530000 2.375000 ;
      RECT 7.710000  2.255000 8.040000 2.635000 ;
      RECT 7.815000  0.465000 8.135000 0.820000 ;
      RECT 7.815000  0.820000 8.140000 0.995000 ;
      RECT 7.815000  0.995000 8.730000 1.295000 ;
      RECT 7.990000  1.295000 8.730000 1.325000 ;
      RECT 7.990000  1.325000 8.160000 1.915000 ;
      RECT 8.380000  0.085000 8.685000 0.545000 ;
      RECT 8.380000  1.495000 8.685000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.105000 0.780000 1.275000 ;
      RECT 1.015000  1.785000 1.185000 1.955000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  1.105000 2.615000 1.275000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  1.785000 3.075000 1.955000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.025000  1.105000 6.195000 1.275000 ;
      RECT 6.025000  1.785000 6.195000 1.955000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.075000 0.840000 1.120000 ;
      RECT 0.550000 1.120000 6.255000 1.260000 ;
      RECT 0.550000 1.260000 0.840000 1.305000 ;
      RECT 0.955000 1.755000 1.245000 1.800000 ;
      RECT 0.955000 1.800000 6.255000 1.940000 ;
      RECT 0.955000 1.940000 1.245000 1.985000 ;
      RECT 2.385000 1.075000 2.675000 1.120000 ;
      RECT 2.385000 1.260000 2.675000 1.305000 ;
      RECT 2.845000 1.755000 3.135000 1.800000 ;
      RECT 2.845000 1.940000 3.135000 1.985000 ;
      RECT 5.965000 1.075000 6.255000 1.120000 ;
      RECT 5.965000 1.260000 6.255000 1.305000 ;
      RECT 5.965000 1.755000 6.255000 1.800000 ;
      RECT 5.965000 1.940000 6.255000 1.985000 ;
  END
END sky130_fd_sc_hd__dfrtp_1
MACRO sky130_fd_sc_hd__dfrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.665000 1.680000 2.450000 ;
        RECT 1.415000 0.615000 1.875000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.855000 0.265000 9.105000 0.795000 ;
        RECT 8.855000 1.445000 9.105000 2.325000 ;
        RECT 8.900000 0.795000 9.105000 1.445000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.765000 4.595000 1.015000 ;
      LAYER mcon ;
        RECT 4.165000 0.765000 4.335000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105000 1.035000 7.645000 1.405000 ;
        RECT 7.405000 0.635000 7.645000 1.035000 ;
      LAYER mcon ;
        RECT 7.105000 1.080000 7.275000 1.250000 ;
        RECT 7.405000 0.765000 7.575000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745000 0.735000 4.395000 0.780000 ;
        RECT 3.745000 0.780000 7.635000 0.920000 ;
        RECT 3.745000 0.920000 4.395000 0.965000 ;
        RECT 7.045000 0.920000 7.635000 0.965000 ;
        RECT 7.045000 0.965000 7.335000 1.280000 ;
        RECT 7.345000 0.735000 7.635000 0.780000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.090000  0.345000 0.345000 0.635000 ;
      RECT 0.090000  0.635000 0.840000 0.805000 ;
      RECT 0.090000  1.795000 0.840000 1.965000 ;
      RECT 0.090000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 2.465000 ;
      RECT 1.545000  0.085000 1.875000 0.445000 ;
      RECT 1.850000  2.175000 2.100000 2.635000 ;
      RECT 2.045000  0.305000 2.540000 0.475000 ;
      RECT 2.045000  0.475000 2.215000 1.835000 ;
      RECT 2.045000  1.835000 2.440000 2.005000 ;
      RECT 2.270000  2.005000 2.440000 2.135000 ;
      RECT 2.270000  2.135000 2.520000 2.465000 ;
      RECT 2.385000  0.765000 2.735000 1.385000 ;
      RECT 2.610000  1.575000 3.075000 1.965000 ;
      RECT 2.735000  2.135000 3.415000 2.465000 ;
      RECT 2.745000  0.305000 3.600000 0.475000 ;
      RECT 2.905000  0.765000 3.260000 0.985000 ;
      RECT 2.905000  0.985000 3.075000 1.575000 ;
      RECT 3.245000  1.185000 4.935000 1.355000 ;
      RECT 3.245000  1.355000 3.415000 2.135000 ;
      RECT 3.430000  0.475000 3.600000 1.185000 ;
      RECT 3.585000  1.865000 4.660000 2.035000 ;
      RECT 3.585000  2.035000 3.755000 2.375000 ;
      RECT 3.775000  1.525000 5.275000 1.695000 ;
      RECT 3.990000  2.205000 4.320000 2.635000 ;
      RECT 4.475000  0.085000 4.805000 0.545000 ;
      RECT 4.490000  2.035000 4.660000 2.375000 ;
      RECT 4.765000  1.005000 4.935000 1.185000 ;
      RECT 4.955000  2.175000 5.325000 2.635000 ;
      RECT 5.015000  0.275000 5.365000 0.445000 ;
      RECT 5.015000  0.445000 5.275000 0.835000 ;
      RECT 5.105000  0.835000 5.275000 1.525000 ;
      RECT 5.105000  1.695000 5.275000 1.835000 ;
      RECT 5.105000  1.835000 5.665000 2.005000 ;
      RECT 5.465000  0.705000 5.675000 1.495000 ;
      RECT 5.465000  1.495000 6.140000 1.655000 ;
      RECT 5.465000  1.655000 6.430000 1.665000 ;
      RECT 5.495000  2.005000 5.665000 2.465000 ;
      RECT 5.585000  0.255000 6.535000 0.535000 ;
      RECT 5.845000  0.705000 6.195000 1.325000 ;
      RECT 5.900000  2.125000 6.770000 2.465000 ;
      RECT 5.970000  1.665000 6.430000 1.955000 ;
      RECT 6.365000  0.535000 6.535000 1.315000 ;
      RECT 6.365000  1.315000 6.770000 1.485000 ;
      RECT 6.600000  1.485000 6.770000 1.575000 ;
      RECT 6.600000  1.575000 7.820000 1.745000 ;
      RECT 6.600000  1.745000 6.770000 2.125000 ;
      RECT 6.705000  0.085000 6.895000 0.525000 ;
      RECT 6.705000  0.695000 7.235000 0.865000 ;
      RECT 6.705000  0.865000 6.925000 1.145000 ;
      RECT 6.940000  2.175000 7.190000 2.635000 ;
      RECT 7.065000  0.295000 8.135000 0.465000 ;
      RECT 7.065000  0.465000 7.235000 0.695000 ;
      RECT 7.360000  1.915000 8.160000 2.085000 ;
      RECT 7.360000  2.085000 7.530000 2.375000 ;
      RECT 7.710000  2.255000 8.040000 2.635000 ;
      RECT 7.815000  0.465000 8.135000 0.820000 ;
      RECT 7.815000  0.820000 8.140000 0.995000 ;
      RECT 7.815000  0.995000 8.730000 1.295000 ;
      RECT 7.990000  1.295000 8.730000 1.325000 ;
      RECT 7.990000  1.325000 8.160000 1.915000 ;
      RECT 8.380000  0.085000 8.685000 0.545000 ;
      RECT 8.380000  1.495000 8.685000 2.635000 ;
      RECT 9.275000  0.085000 9.525000 0.840000 ;
      RECT 9.275000  1.495000 9.525000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.105000 0.780000 1.275000 ;
      RECT 1.015000  1.785000 1.185000 1.955000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  1.105000 2.615000 1.275000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  1.785000 3.075000 1.955000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.025000  1.105000 6.195000 1.275000 ;
      RECT 6.025000  1.785000 6.195000 1.955000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.075000 0.840000 1.120000 ;
      RECT 0.550000 1.120000 6.255000 1.260000 ;
      RECT 0.550000 1.260000 0.840000 1.305000 ;
      RECT 0.955000 1.755000 1.245000 1.800000 ;
      RECT 0.955000 1.800000 6.255000 1.940000 ;
      RECT 0.955000 1.940000 1.245000 1.985000 ;
      RECT 2.385000 1.075000 2.675000 1.120000 ;
      RECT 2.385000 1.260000 2.675000 1.305000 ;
      RECT 2.845000 1.755000 3.135000 1.800000 ;
      RECT 2.845000 1.940000 3.135000 1.985000 ;
      RECT 5.965000 1.075000 6.255000 1.120000 ;
      RECT 5.965000 1.260000 6.255000 1.305000 ;
      RECT 5.965000 1.755000 6.255000 1.800000 ;
      RECT 5.965000 1.940000 6.255000 1.985000 ;
  END
END sky130_fd_sc_hd__dfrtp_2
MACRO sky130_fd_sc_hd__dfrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.58000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.665000 1.680000 2.450000 ;
        RECT 1.415000 0.615000 1.875000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  8.675000 0.255000  9.005000 0.735000 ;
        RECT  8.675000 0.735000 10.440000 0.905000 ;
        RECT  8.715000 1.455000 10.440000 1.625000 ;
        RECT  8.715000 1.625000  9.005000 2.465000 ;
        RECT  9.515000 0.255000  9.845000 0.735000 ;
        RECT  9.555000 1.625000  9.805000 2.465000 ;
        RECT 10.030000 0.905000 10.440000 1.455000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.765000 4.595000 1.015000 ;
      LAYER mcon ;
        RECT 4.165000 0.765000 4.335000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105000 1.035000 7.645000 1.405000 ;
        RECT 7.405000 0.635000 7.645000 1.035000 ;
      LAYER mcon ;
        RECT 7.105000 1.080000 7.275000 1.250000 ;
        RECT 7.405000 0.765000 7.575000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745000 0.735000 4.395000 0.780000 ;
        RECT 3.745000 0.780000 7.635000 0.920000 ;
        RECT 3.745000 0.920000 4.395000 0.965000 ;
        RECT 7.045000 0.920000 7.635000 0.965000 ;
        RECT 7.045000 0.965000 7.335000 1.280000 ;
        RECT 7.345000 0.735000 7.635000 0.780000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.770000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.580000 0.085000 ;
      RECT  0.000000  2.635000 10.580000 2.805000 ;
      RECT  0.090000  0.345000  0.345000 0.635000 ;
      RECT  0.090000  0.635000  0.840000 0.805000 ;
      RECT  0.090000  1.795000  0.840000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.610000  0.805000  0.840000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.545000  0.085000  1.875000 0.445000 ;
      RECT  1.850000  2.175000  2.100000 2.635000 ;
      RECT  2.045000  0.305000  2.540000 0.475000 ;
      RECT  2.045000  0.475000  2.215000 1.835000 ;
      RECT  2.045000  1.835000  2.440000 2.005000 ;
      RECT  2.270000  2.005000  2.440000 2.135000 ;
      RECT  2.270000  2.135000  2.520000 2.465000 ;
      RECT  2.385000  0.765000  2.735000 1.385000 ;
      RECT  2.610000  1.575000  3.075000 1.965000 ;
      RECT  2.735000  2.135000  3.415000 2.465000 ;
      RECT  2.745000  0.305000  3.600000 0.475000 ;
      RECT  2.905000  0.765000  3.260000 0.985000 ;
      RECT  2.905000  0.985000  3.075000 1.575000 ;
      RECT  3.245000  1.185000  4.935000 1.355000 ;
      RECT  3.245000  1.355000  3.415000 2.135000 ;
      RECT  3.430000  0.475000  3.600000 1.185000 ;
      RECT  3.585000  1.865000  4.660000 2.035000 ;
      RECT  3.585000  2.035000  3.755000 2.375000 ;
      RECT  3.775000  1.525000  5.275000 1.695000 ;
      RECT  3.990000  2.205000  4.320000 2.635000 ;
      RECT  4.475000  0.085000  4.805000 0.545000 ;
      RECT  4.490000  2.035000  4.660000 2.375000 ;
      RECT  4.765000  1.005000  4.935000 1.185000 ;
      RECT  4.955000  2.175000  5.325000 2.635000 ;
      RECT  5.015000  0.275000  5.365000 0.445000 ;
      RECT  5.015000  0.445000  5.275000 0.835000 ;
      RECT  5.105000  0.835000  5.275000 1.525000 ;
      RECT  5.105000  1.695000  5.275000 1.835000 ;
      RECT  5.105000  1.835000  5.665000 2.005000 ;
      RECT  5.465000  0.705000  5.675000 1.495000 ;
      RECT  5.465000  1.495000  6.140000 1.655000 ;
      RECT  5.465000  1.655000  6.430000 1.665000 ;
      RECT  5.495000  2.005000  5.665000 2.465000 ;
      RECT  5.585000  0.255000  6.535000 0.535000 ;
      RECT  5.845000  0.705000  6.195000 1.325000 ;
      RECT  5.900000  2.125000  6.770000 2.465000 ;
      RECT  5.970000  1.665000  6.430000 1.955000 ;
      RECT  6.365000  0.535000  6.535000 1.315000 ;
      RECT  6.365000  1.315000  6.770000 1.485000 ;
      RECT  6.600000  1.485000  6.770000 1.575000 ;
      RECT  6.600000  1.575000  7.820000 1.745000 ;
      RECT  6.600000  1.745000  6.770000 2.125000 ;
      RECT  6.705000  0.085000  6.895000 0.525000 ;
      RECT  6.705000  0.695000  7.235000 0.865000 ;
      RECT  6.705000  0.865000  6.925000 1.145000 ;
      RECT  6.940000  2.175000  7.190000 2.635000 ;
      RECT  7.065000  0.295000  8.135000 0.465000 ;
      RECT  7.065000  0.465000  7.235000 0.695000 ;
      RECT  7.360000  1.915000  8.160000 2.085000 ;
      RECT  7.360000  2.085000  7.530000 2.375000 ;
      RECT  7.710000  2.255000  8.040000 2.635000 ;
      RECT  7.815000  0.465000  8.135000 0.820000 ;
      RECT  7.815000  0.820000  8.140000 1.075000 ;
      RECT  7.815000  1.075000  9.845000 1.285000 ;
      RECT  7.815000  1.285000  8.160000 1.295000 ;
      RECT  7.990000  1.295000  8.160000 1.915000 ;
      RECT  8.335000  0.085000  8.505000 0.895000 ;
      RECT  8.335000  1.575000  8.505000 2.635000 ;
      RECT  9.175000  0.085000  9.345000 0.555000 ;
      RECT  9.175000  1.795000  9.345000 2.635000 ;
      RECT 10.015000  0.085000 10.185000 0.555000 ;
      RECT 10.015000  1.795000 10.185000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.610000  1.105000  0.780000 1.275000 ;
      RECT  1.015000  1.785000  1.185000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  1.105000  2.615000 1.275000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  1.785000  3.075000 1.955000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.025000  1.105000  6.195000 1.275000 ;
      RECT  6.025000  1.785000  6.195000 1.955000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.075000 0.840000 1.120000 ;
      RECT 0.550000 1.120000 6.255000 1.260000 ;
      RECT 0.550000 1.260000 0.840000 1.305000 ;
      RECT 0.955000 1.755000 1.245000 1.800000 ;
      RECT 0.955000 1.800000 6.255000 1.940000 ;
      RECT 0.955000 1.940000 1.245000 1.985000 ;
      RECT 2.385000 1.075000 2.675000 1.120000 ;
      RECT 2.385000 1.260000 2.675000 1.305000 ;
      RECT 2.845000 1.755000 3.135000 1.800000 ;
      RECT 2.845000 1.940000 3.135000 1.985000 ;
      RECT 5.965000 1.075000 6.255000 1.120000 ;
      RECT 5.965000 1.260000 6.255000 1.305000 ;
      RECT 5.965000 1.755000 6.255000 1.800000 ;
      RECT 5.965000 1.940000 6.255000 1.985000 ;
  END
END sky130_fd_sc_hd__dfrtp_4
MACRO sky130_fd_sc_hd__dfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfsbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.58000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.770000 1.005000 2.180000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.865000 0.255000 10.125000 0.825000 ;
        RECT 9.865000 1.445000 10.125000 2.465000 ;
        RECT 9.910000 0.825000 10.125000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.370000 0.255000 8.700000 2.465000 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.610000 0.735000 4.020000 1.065000 ;
      LAYER mcon ;
        RECT 3.825000 0.765000 3.995000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.660000 0.735000 7.320000 1.005000 ;
        RECT 6.660000 1.005000 6.990000 1.065000 ;
      LAYER mcon ;
        RECT 7.045000 0.765000 7.215000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765000 0.735000 4.055000 0.780000 ;
        RECT 3.765000 0.780000 7.275000 0.920000 ;
        RECT 3.765000 0.920000 4.055000 0.965000 ;
        RECT 6.985000 0.735000 7.275000 0.780000 ;
        RECT 6.985000 0.920000 7.275000 0.965000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.770000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.580000 0.085000 ;
      RECT 0.000000  2.635000 10.580000 2.805000 ;
      RECT 0.175000  0.345000  0.345000 0.635000 ;
      RECT 0.175000  0.635000  0.840000 0.805000 ;
      RECT 0.175000  1.795000  0.840000 1.965000 ;
      RECT 0.175000  1.965000  0.345000 2.465000 ;
      RECT 0.515000  0.085000  0.845000 0.465000 ;
      RECT 0.515000  2.135000  0.845000 2.635000 ;
      RECT 0.610000  0.805000  0.840000 1.795000 ;
      RECT 1.015000  0.345000  1.240000 2.465000 ;
      RECT 1.430000  0.635000  2.125000 0.825000 ;
      RECT 1.430000  0.825000  1.600000 1.795000 ;
      RECT 1.430000  1.795000  2.125000 1.965000 ;
      RECT 1.455000  0.085000  1.785000 0.465000 ;
      RECT 1.455000  2.135000  1.785000 2.635000 ;
      RECT 1.955000  0.305000  2.125000 0.635000 ;
      RECT 1.955000  1.965000  2.125000 2.465000 ;
      RECT 2.350000  0.705000  2.570000 1.575000 ;
      RECT 2.350000  1.575000  2.850000 1.955000 ;
      RECT 2.360000  2.250000  3.190000 2.420000 ;
      RECT 2.425000  0.265000  3.440000 0.465000 ;
      RECT 2.750000  0.645000  3.100000 1.015000 ;
      RECT 3.020000  1.195000  3.440000 1.235000 ;
      RECT 3.020000  1.235000  4.370000 1.405000 ;
      RECT 3.020000  1.405000  3.190000 2.250000 ;
      RECT 3.270000  0.465000  3.440000 1.195000 ;
      RECT 3.360000  1.575000  3.610000 1.835000 ;
      RECT 3.360000  1.835000  4.710000 2.085000 ;
      RECT 3.430000  2.255000  3.810000 2.635000 ;
      RECT 3.610000  0.085000  4.020000 0.525000 ;
      RECT 3.990000  2.085000  4.160000 2.375000 ;
      RECT 4.120000  1.405000  4.370000 1.565000 ;
      RECT 4.310000  0.295000  4.560000 0.725000 ;
      RECT 4.310000  0.725000  4.710000 1.065000 ;
      RECT 4.330000  2.255000  4.660000 2.635000 ;
      RECT 4.540000  1.065000  4.710000 1.835000 ;
      RECT 4.740000  0.085000  5.080000 0.545000 ;
      RECT 4.900000  0.725000  6.150000 0.895000 ;
      RECT 4.900000  0.895000  5.070000 1.655000 ;
      RECT 4.900000  1.655000  5.400000 1.965000 ;
      RECT 5.110000  2.165000  5.760000 2.415000 ;
      RECT 5.240000  1.065000  5.420000 1.475000 ;
      RECT 5.590000  1.235000  7.470000 1.405000 ;
      RECT 5.590000  1.405000  5.760000 1.915000 ;
      RECT 5.590000  1.915000  6.780000 2.085000 ;
      RECT 5.590000  2.085000  5.760000 2.165000 ;
      RECT 5.640000  0.305000  6.490000 0.475000 ;
      RECT 5.820000  0.895000  6.150000 1.015000 ;
      RECT 5.930000  1.575000  7.830000 1.745000 ;
      RECT 5.930000  2.255000  6.340000 2.635000 ;
      RECT 6.320000  0.475000  6.490000 1.235000 ;
      RECT 6.540000  2.085000  6.780000 2.375000 ;
      RECT 6.670000  0.085000  7.330000 0.565000 ;
      RECT 7.010000  1.945000  7.340000 2.635000 ;
      RECT 7.140000  1.175000  7.470000 1.235000 ;
      RECT 7.510000  0.350000  7.830000 0.680000 ;
      RECT 7.510000  1.745000  7.830000 1.765000 ;
      RECT 7.510000  1.765000  7.680000 2.375000 ;
      RECT 7.640000  0.680000  7.830000 1.575000 ;
      RECT 8.020000  0.085000  8.200000 0.905000 ;
      RECT 8.020000  1.480000  8.200000 2.635000 ;
      RECT 8.890000  0.255000  9.220000 0.995000 ;
      RECT 8.890000  0.995000  9.740000 1.325000 ;
      RECT 8.890000  1.325000  9.220000 2.465000 ;
      RECT 9.445000  0.085000  9.615000 0.585000 ;
      RECT 9.445000  1.825000  9.615000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.645000  1.785000  0.815000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  0.765000  1.235000 0.935000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  1.785000  2.615000 1.955000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  0.765000  3.075000 0.935000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.245000  1.105000  5.415000 1.275000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
    LAYER met1 ;
      RECT 0.585000 1.755000 0.875000 1.800000 ;
      RECT 0.585000 1.800000 5.435000 1.940000 ;
      RECT 0.585000 1.940000 0.875000 1.985000 ;
      RECT 1.005000 0.735000 1.295000 0.780000 ;
      RECT 1.005000 0.780000 3.135000 0.920000 ;
      RECT 1.005000 0.920000 1.295000 0.965000 ;
      RECT 2.385000 1.755000 2.675000 1.800000 ;
      RECT 2.385000 1.940000 2.675000 1.985000 ;
      RECT 2.845000 0.735000 3.135000 0.780000 ;
      RECT 2.845000 0.920000 3.135000 0.965000 ;
      RECT 2.920000 0.965000 3.135000 1.120000 ;
      RECT 2.920000 1.120000 5.475000 1.260000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 5.185000 1.075000 5.475000 1.120000 ;
      RECT 5.185000 1.260000 5.475000 1.305000 ;
  END
END sky130_fd_sc_hd__dfsbp_1
MACRO sky130_fd_sc_hd__dfsbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfsbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.770000 1.005000 2.180000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.150000 1.495000 10.915000 1.665000 ;
        RECT 10.150000 1.665000 10.480000 2.465000 ;
        RECT 10.230000 0.255000 10.480000 0.720000 ;
        RECT 10.230000 0.720000 10.915000 0.825000 ;
        RECT 10.345000 0.825000 10.915000 0.845000 ;
        RECT 10.360000 0.845000 10.915000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.370000 0.255000 8.700000 2.465000 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.610000 0.735000 4.020000 1.065000 ;
      LAYER mcon ;
        RECT 3.825000 0.765000 3.995000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.660000 0.735000 7.320000 1.005000 ;
        RECT 6.660000 1.005000 6.990000 1.065000 ;
      LAYER mcon ;
        RECT 7.045000 0.765000 7.215000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765000 0.735000 4.055000 0.780000 ;
        RECT 3.765000 0.780000 7.275000 0.920000 ;
        RECT 3.765000 0.920000 4.055000 0.965000 ;
        RECT 6.985000 0.735000 7.275000 0.780000 ;
        RECT 6.985000 0.920000 7.275000 0.965000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.840000 0.805000 ;
      RECT  0.175000  1.795000  0.840000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.610000  0.805000  0.840000 1.795000 ;
      RECT  1.015000  0.345000  1.240000 2.465000 ;
      RECT  1.430000  0.635000  2.125000 0.825000 ;
      RECT  1.430000  0.825000  1.600000 1.795000 ;
      RECT  1.430000  1.795000  2.125000 1.965000 ;
      RECT  1.455000  0.085000  1.785000 0.465000 ;
      RECT  1.455000  2.135000  1.785000 2.635000 ;
      RECT  1.955000  0.305000  2.125000 0.635000 ;
      RECT  1.955000  1.965000  2.125000 2.465000 ;
      RECT  2.350000  0.705000  2.570000 1.575000 ;
      RECT  2.350000  1.575000  2.850000 1.955000 ;
      RECT  2.360000  2.250000  3.190000 2.420000 ;
      RECT  2.425000  0.265000  3.440000 0.465000 ;
      RECT  2.750000  0.645000  3.100000 1.015000 ;
      RECT  3.020000  1.195000  3.440000 1.235000 ;
      RECT  3.020000  1.235000  4.370000 1.405000 ;
      RECT  3.020000  1.405000  3.190000 2.250000 ;
      RECT  3.270000  0.465000  3.440000 1.195000 ;
      RECT  3.360000  1.575000  3.610000 1.835000 ;
      RECT  3.360000  1.835000  4.710000 2.085000 ;
      RECT  3.430000  2.255000  3.810000 2.635000 ;
      RECT  3.610000  0.085000  4.020000 0.525000 ;
      RECT  3.990000  2.085000  4.160000 2.375000 ;
      RECT  4.120000  1.405000  4.370000 1.565000 ;
      RECT  4.310000  0.295000  4.560000 0.725000 ;
      RECT  4.310000  0.725000  4.710000 1.065000 ;
      RECT  4.330000  2.255000  4.660000 2.635000 ;
      RECT  4.540000  1.065000  4.710000 1.835000 ;
      RECT  4.740000  0.085000  5.080000 0.545000 ;
      RECT  4.900000  0.725000  6.150000 0.895000 ;
      RECT  4.900000  0.895000  5.070000 1.655000 ;
      RECT  4.900000  1.655000  5.400000 1.965000 ;
      RECT  5.110000  2.165000  5.760000 2.415000 ;
      RECT  5.240000  1.065000  5.420000 1.475000 ;
      RECT  5.590000  1.235000  7.470000 1.405000 ;
      RECT  5.590000  1.405000  5.760000 1.915000 ;
      RECT  5.590000  1.915000  6.780000 2.085000 ;
      RECT  5.590000  2.085000  5.760000 2.165000 ;
      RECT  5.640000  0.305000  6.490000 0.475000 ;
      RECT  5.820000  0.895000  6.150000 1.015000 ;
      RECT  5.930000  1.575000  7.830000 1.745000 ;
      RECT  5.930000  2.255000  6.340000 2.635000 ;
      RECT  6.320000  0.475000  6.490000 1.235000 ;
      RECT  6.540000  2.085000  6.780000 2.375000 ;
      RECT  6.670000  0.085000  7.330000 0.565000 ;
      RECT  7.010000  1.945000  7.340000 2.635000 ;
      RECT  7.140000  1.175000  7.470000 1.235000 ;
      RECT  7.510000  0.350000  7.830000 0.680000 ;
      RECT  7.510000  1.745000  7.830000 1.765000 ;
      RECT  7.510000  1.765000  7.680000 2.375000 ;
      RECT  7.640000  0.680000  7.830000 1.575000 ;
      RECT  8.020000  0.085000  8.200000 0.905000 ;
      RECT  8.020000  1.480000  8.200000 2.635000 ;
      RECT  8.870000  0.085000  9.120000 0.905000 ;
      RECT  8.870000  1.480000  9.120000 2.635000 ;
      RECT  9.310000  0.255000  9.560000 0.995000 ;
      RECT  9.310000  0.995000 10.190000 1.325000 ;
      RECT  9.310000  1.325000  9.640000 2.465000 ;
      RECT  9.730000  0.085000 10.060000 0.825000 ;
      RECT  9.810000  1.495000  9.980000 2.635000 ;
      RECT 10.650000  0.085000 10.915000 0.550000 ;
      RECT 10.650000  1.835000 10.915000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.645000  1.785000  0.815000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  0.765000  1.235000 0.935000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  1.785000  2.615000 1.955000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  0.765000  3.075000 0.935000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.245000  1.105000  5.415000 1.275000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 0.585000 1.755000 0.875000 1.800000 ;
      RECT 0.585000 1.800000 5.435000 1.940000 ;
      RECT 0.585000 1.940000 0.875000 1.985000 ;
      RECT 1.005000 0.735000 1.295000 0.780000 ;
      RECT 1.005000 0.780000 3.135000 0.920000 ;
      RECT 1.005000 0.920000 1.295000 0.965000 ;
      RECT 2.385000 1.755000 2.675000 1.800000 ;
      RECT 2.385000 1.940000 2.675000 1.985000 ;
      RECT 2.845000 0.735000 3.135000 0.780000 ;
      RECT 2.845000 0.920000 3.135000 0.965000 ;
      RECT 2.920000 0.965000 3.135000 1.120000 ;
      RECT 2.920000 1.120000 5.475000 1.260000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 5.185000 1.075000 5.475000 1.120000 ;
      RECT 5.185000 1.260000 5.475000 1.305000 ;
  END
END sky130_fd_sc_hd__dfsbp_2
MACRO sky130_fd_sc_hd__dfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfstp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.770000 1.005000 2.180000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.945000 0.265000 9.200000 0.795000 ;
        RECT 8.945000 1.655000 9.200000 2.325000 ;
        RECT 9.020000 0.795000 9.200000 1.655000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.610000 0.735000 4.020000 1.065000 ;
      LAYER mcon ;
        RECT 3.850000 0.765000 4.020000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.680000 0.735000 7.340000 1.005000 ;
        RECT 6.680000 1.005000 7.010000 1.065000 ;
      LAYER mcon ;
        RECT 7.110000 0.765000 7.280000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.790000 0.735000 4.080000 0.780000 ;
        RECT 3.790000 0.780000 7.340000 0.920000 ;
        RECT 3.790000 0.920000 4.080000 0.965000 ;
        RECT 7.050000 0.735000 7.340000 0.780000 ;
        RECT 7.050000 0.920000 7.340000 0.965000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.840000 0.805000 ;
      RECT 0.175000  1.795000 0.840000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.240000 2.465000 ;
      RECT 1.430000  0.635000 2.125000 0.825000 ;
      RECT 1.430000  0.825000 1.600000 1.795000 ;
      RECT 1.430000  1.795000 2.125000 1.965000 ;
      RECT 1.455000  0.085000 1.785000 0.465000 ;
      RECT 1.455000  2.135000 1.785000 2.635000 ;
      RECT 1.955000  0.305000 2.125000 0.635000 ;
      RECT 1.955000  1.965000 2.125000 2.465000 ;
      RECT 2.350000  0.705000 2.570000 1.575000 ;
      RECT 2.350000  1.575000 2.850000 1.955000 ;
      RECT 2.360000  2.250000 3.190000 2.420000 ;
      RECT 2.425000  0.265000 3.440000 0.465000 ;
      RECT 2.750000  0.645000 3.100000 1.015000 ;
      RECT 3.020000  1.195000 3.440000 1.235000 ;
      RECT 3.020000  1.235000 4.370000 1.405000 ;
      RECT 3.020000  1.405000 3.190000 2.250000 ;
      RECT 3.270000  0.465000 3.440000 1.195000 ;
      RECT 3.360000  1.575000 3.610000 1.835000 ;
      RECT 3.360000  1.835000 4.730000 2.085000 ;
      RECT 3.430000  2.255000 3.810000 2.635000 ;
      RECT 3.610000  0.085000 4.020000 0.525000 ;
      RECT 3.990000  2.085000 4.160000 2.375000 ;
      RECT 4.120000  1.405000 4.370000 1.565000 ;
      RECT 4.310000  0.295000 4.560000 0.725000 ;
      RECT 4.310000  0.725000 4.730000 1.065000 ;
      RECT 4.330000  2.255000 4.660000 2.635000 ;
      RECT 4.540000  1.065000 4.730000 1.835000 ;
      RECT 4.760000  0.085000 5.080000 0.545000 ;
      RECT 4.900000  0.725000 6.150000 0.895000 ;
      RECT 4.900000  0.895000 5.070000 1.655000 ;
      RECT 4.900000  1.655000 5.420000 1.965000 ;
      RECT 5.130000  2.165000 5.760000 2.415000 ;
      RECT 5.240000  1.065000 5.420000 1.475000 ;
      RECT 5.590000  1.235000 7.490000 1.405000 ;
      RECT 5.590000  1.405000 5.760000 1.915000 ;
      RECT 5.590000  1.915000 6.800000 2.085000 ;
      RECT 5.590000  2.085000 5.760000 2.165000 ;
      RECT 5.640000  0.305000 6.490000 0.475000 ;
      RECT 5.820000  0.895000 6.150000 1.015000 ;
      RECT 5.930000  1.575000 7.850000 1.745000 ;
      RECT 5.940000  2.255000 6.360000 2.635000 ;
      RECT 6.320000  0.475000 6.490000 1.235000 ;
      RECT 6.560000  2.085000 6.800000 2.375000 ;
      RECT 6.690000  0.085000 7.350000 0.565000 ;
      RECT 7.030000  1.945000 7.360000 2.635000 ;
      RECT 7.160000  1.175000 7.490000 1.235000 ;
      RECT 7.530000  0.350000 7.850000 0.680000 ;
      RECT 7.530000  1.745000 7.850000 1.765000 ;
      RECT 7.530000  1.765000 7.700000 2.375000 ;
      RECT 7.660000  0.680000 7.850000 1.575000 ;
      RECT 7.970000  1.915000 8.300000 2.425000 ;
      RECT 8.050000  0.345000 8.300000 0.995000 ;
      RECT 8.050000  0.995000 8.850000 1.325000 ;
      RECT 8.050000  1.325000 8.300000 1.915000 ;
      RECT 8.480000  0.085000 8.765000 0.545000 ;
      RECT 8.480000  1.835000 8.765000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.785000 0.780000 1.955000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  0.765000 1.240000 0.935000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.785000 2.640000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  0.765000 3.100000 0.935000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.250000  1.105000 5.420000 1.275000 ;
      RECT 5.250000  1.785000 5.420000 1.955000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.755000 0.840000 1.800000 ;
      RECT 0.550000 1.800000 5.480000 1.940000 ;
      RECT 0.550000 1.940000 0.840000 1.985000 ;
      RECT 1.010000 0.735000 1.300000 0.780000 ;
      RECT 1.010000 0.780000 3.160000 0.920000 ;
      RECT 1.010000 0.920000 1.300000 0.965000 ;
      RECT 2.410000 1.755000 2.700000 1.800000 ;
      RECT 2.410000 1.940000 2.700000 1.985000 ;
      RECT 2.870000 0.735000 3.160000 0.780000 ;
      RECT 2.870000 0.920000 3.160000 0.965000 ;
      RECT 2.945000 0.965000 3.160000 1.120000 ;
      RECT 2.945000 1.120000 5.480000 1.260000 ;
      RECT 5.190000 1.075000 5.480000 1.120000 ;
      RECT 5.190000 1.260000 5.480000 1.305000 ;
      RECT 5.190000 1.755000 5.480000 1.800000 ;
      RECT 5.190000 1.940000 5.480000 1.985000 ;
  END
END sky130_fd_sc_hd__dfstp_1
MACRO sky130_fd_sc_hd__dfstp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfstp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.770000 1.005000 2.180000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.810000 1.495000 9.575000 1.615000 ;
        RECT 8.810000 1.615000 9.140000 2.460000 ;
        RECT 8.890000 0.265000 9.135000 0.765000 ;
        RECT 8.890000 0.765000 9.575000 0.825000 ;
        RECT 8.975000 0.825000 9.575000 0.855000 ;
        RECT 8.975000 1.445000 9.575000 1.495000 ;
        RECT 8.990000 0.855000 9.575000 0.895000 ;
        RECT 9.020000 0.895000 9.575000 1.445000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.610000 0.735000 4.020000 1.065000 ;
      LAYER mcon ;
        RECT 3.825000 0.765000 3.995000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.660000 0.735000 7.340000 1.005000 ;
        RECT 6.660000 1.005000 7.010000 1.065000 ;
      LAYER mcon ;
        RECT 7.045000 0.765000 7.215000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765000 0.735000 4.055000 0.780000 ;
        RECT 3.765000 0.780000 7.275000 0.920000 ;
        RECT 3.765000 0.920000 4.055000 0.965000 ;
        RECT 6.985000 0.735000 7.275000 0.780000 ;
        RECT 6.985000 0.920000 7.275000 0.965000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.435000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.635000 ;
      RECT 0.085000  0.635000 0.835000 0.805000 ;
      RECT 0.085000  1.795000 0.835000 1.965000 ;
      RECT 0.085000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.605000  0.805000 0.835000 1.795000 ;
      RECT 1.005000  0.565000 1.235000 2.045000 ;
      RECT 1.015000  0.345000 1.235000 0.565000 ;
      RECT 1.015000  2.045000 1.235000 2.465000 ;
      RECT 1.430000  0.635000 2.125000 0.825000 ;
      RECT 1.430000  0.825000 1.600000 1.795000 ;
      RECT 1.430000  1.795000 2.125000 1.965000 ;
      RECT 1.455000  0.085000 1.785000 0.465000 ;
      RECT 1.455000  2.135000 1.785000 2.635000 ;
      RECT 1.955000  0.305000 2.125000 0.635000 ;
      RECT 1.955000  1.965000 2.125000 2.465000 ;
      RECT 2.350000  0.705000 2.570000 1.575000 ;
      RECT 2.350000  1.575000 2.850000 1.955000 ;
      RECT 2.360000  2.250000 3.190000 2.420000 ;
      RECT 2.425000  0.265000 3.440000 0.465000 ;
      RECT 2.750000  0.645000 3.100000 1.015000 ;
      RECT 3.020000  1.195000 3.440000 1.235000 ;
      RECT 3.020000  1.235000 4.370000 1.405000 ;
      RECT 3.020000  1.405000 3.190000 2.250000 ;
      RECT 3.270000  0.465000 3.440000 1.195000 ;
      RECT 3.360000  1.575000 3.610000 1.835000 ;
      RECT 3.360000  1.835000 4.710000 2.085000 ;
      RECT 3.430000  2.255000 3.810000 2.635000 ;
      RECT 3.610000  0.085000 4.020000 0.525000 ;
      RECT 3.990000  2.085000 4.160000 2.375000 ;
      RECT 4.120000  1.405000 4.370000 1.565000 ;
      RECT 4.310000  0.295000 4.560000 0.725000 ;
      RECT 4.310000  0.725000 4.710000 1.065000 ;
      RECT 4.330000  2.255000 4.660000 2.635000 ;
      RECT 4.540000  1.065000 4.710000 1.835000 ;
      RECT 4.760000  0.085000 5.080000 0.545000 ;
      RECT 4.880000  0.725000 6.150000 0.895000 ;
      RECT 4.880000  0.895000 5.050000 1.655000 ;
      RECT 4.880000  1.655000 5.400000 1.965000 ;
      RECT 5.110000  2.165000 5.740000 2.415000 ;
      RECT 5.220000  1.065000 5.400000 1.475000 ;
      RECT 5.570000  1.235000 7.490000 1.405000 ;
      RECT 5.570000  1.405000 5.740000 1.915000 ;
      RECT 5.570000  1.915000 6.780000 2.085000 ;
      RECT 5.570000  2.085000 5.740000 2.165000 ;
      RECT 5.640000  0.305000 6.490000 0.475000 ;
      RECT 5.800000  0.895000 6.150000 1.015000 ;
      RECT 5.910000  1.575000 7.880000 1.745000 ;
      RECT 5.920000  2.255000 6.340000 2.635000 ;
      RECT 6.320000  0.475000 6.490000 1.235000 ;
      RECT 6.540000  2.085000 6.780000 2.375000 ;
      RECT 6.690000  0.085000 7.330000 0.565000 ;
      RECT 7.010000  1.945000 7.340000 2.635000 ;
      RECT 7.140000  1.175000 7.490000 1.235000 ;
      RECT 7.510000  1.745000 7.880000 1.765000 ;
      RECT 7.510000  1.765000 7.680000 2.375000 ;
      RECT 7.530000  0.350000 7.880000 0.680000 ;
      RECT 7.690000  0.680000 7.880000 1.575000 ;
      RECT 7.970000  1.915000 8.300000 2.425000 ;
      RECT 8.050000  0.345000 8.220000 0.995000 ;
      RECT 8.050000  0.995000 8.850000 1.325000 ;
      RECT 8.050000  1.325000 8.300000 1.915000 ;
      RECT 8.390000  0.085000 8.720000 0.825000 ;
      RECT 8.470000  1.495000 8.640000 2.635000 ;
      RECT 9.305000  0.085000 9.575000 0.595000 ;
      RECT 9.310000  1.785000 9.575000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  1.785000 0.775000 1.955000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  0.765000 1.235000 0.935000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  1.785000 2.615000 1.955000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  0.765000 3.075000 0.935000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  1.785000 5.375000 1.955000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.225000  1.105000 5.395000 1.275000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 0.545000 1.755000 0.835000 1.800000 ;
      RECT 0.545000 1.800000 5.435000 1.940000 ;
      RECT 0.545000 1.940000 0.835000 1.985000 ;
      RECT 1.005000 0.735000 1.295000 0.780000 ;
      RECT 1.005000 0.780000 3.135000 0.920000 ;
      RECT 1.005000 0.920000 1.295000 0.965000 ;
      RECT 2.385000 1.755000 2.675000 1.800000 ;
      RECT 2.385000 1.940000 2.675000 1.985000 ;
      RECT 2.845000 0.735000 3.135000 0.780000 ;
      RECT 2.845000 0.920000 3.135000 0.965000 ;
      RECT 2.920000 0.965000 3.135000 1.120000 ;
      RECT 2.920000 1.120000 5.455000 1.260000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 5.165000 1.075000 5.455000 1.120000 ;
      RECT 5.165000 1.260000 5.455000 1.305000 ;
  END
END sky130_fd_sc_hd__dfstp_2
MACRO sky130_fd_sc_hd__dfstp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfstp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.770000 1.005000 2.180000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.320000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  8.925000 0.265000  9.170000 0.715000 ;
        RECT  8.925000 0.715000 10.955000 0.885000 ;
        RECT  8.925000 1.470000 10.955000 1.640000 ;
        RECT  8.925000 1.640000  9.170000 2.465000 ;
        RECT  9.765000 0.265000  9.935000 0.715000 ;
        RECT  9.765000 1.640000  9.935000 2.465000 ;
        RECT 10.605000 0.265000 10.955000 0.715000 ;
        RECT 10.605000 1.640000 10.955000 2.465000 ;
        RECT 10.725000 0.885000 10.955000 1.470000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.610000 0.735000 4.020000 1.065000 ;
      LAYER mcon ;
        RECT 3.825000 0.765000 3.995000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.660000 0.735000 7.320000 1.005000 ;
        RECT 6.660000 1.005000 6.990000 1.065000 ;
      LAYER mcon ;
        RECT 7.045000 0.765000 7.215000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765000 0.735000 4.055000 0.780000 ;
        RECT 3.765000 0.780000 7.275000 0.920000 ;
        RECT 3.765000 0.920000 4.055000 0.965000 ;
        RECT 6.985000 0.735000 7.275000 0.780000 ;
        RECT 6.985000 0.920000 7.275000 0.965000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.840000 0.805000 ;
      RECT  0.175000  1.795000  0.840000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.610000  0.805000  0.840000 1.795000 ;
      RECT  1.015000  0.345000  1.240000 2.465000 ;
      RECT  1.430000  0.635000  2.125000 0.825000 ;
      RECT  1.430000  0.825000  1.600000 1.795000 ;
      RECT  1.430000  1.795000  2.125000 1.965000 ;
      RECT  1.455000  0.085000  1.785000 0.465000 ;
      RECT  1.455000  2.135000  1.785000 2.635000 ;
      RECT  1.955000  0.305000  2.125000 0.635000 ;
      RECT  1.955000  1.965000  2.125000 2.465000 ;
      RECT  2.350000  0.705000  2.570000 1.575000 ;
      RECT  2.350000  1.575000  2.850000 1.955000 ;
      RECT  2.360000  2.250000  3.190000 2.420000 ;
      RECT  2.425000  0.265000  3.440000 0.465000 ;
      RECT  2.750000  0.645000  3.100000 1.015000 ;
      RECT  3.020000  1.195000  3.440000 1.235000 ;
      RECT  3.020000  1.235000  4.370000 1.405000 ;
      RECT  3.020000  1.405000  3.190000 2.250000 ;
      RECT  3.270000  0.465000  3.440000 1.195000 ;
      RECT  3.360000  1.575000  3.610000 1.835000 ;
      RECT  3.360000  1.835000  4.710000 2.085000 ;
      RECT  3.430000  2.255000  3.810000 2.635000 ;
      RECT  3.610000  0.085000  4.020000 0.525000 ;
      RECT  3.990000  2.085000  4.160000 2.375000 ;
      RECT  4.120000  1.405000  4.370000 1.565000 ;
      RECT  4.310000  0.295000  4.560000 0.725000 ;
      RECT  4.310000  0.725000  4.710000 1.065000 ;
      RECT  4.330000  2.255000  4.660000 2.635000 ;
      RECT  4.540000  1.065000  4.710000 1.835000 ;
      RECT  4.740000  0.085000  5.080000 0.545000 ;
      RECT  4.880000  0.725000  6.150000 0.895000 ;
      RECT  4.880000  0.895000  5.050000 1.655000 ;
      RECT  4.880000  1.655000  5.400000 1.965000 ;
      RECT  5.110000  2.165000  5.740000 2.415000 ;
      RECT  5.220000  1.065000  5.400000 1.475000 ;
      RECT  5.570000  1.235000  7.470000 1.405000 ;
      RECT  5.570000  1.405000  5.740000 1.915000 ;
      RECT  5.570000  1.915000  6.780000 2.085000 ;
      RECT  5.570000  2.085000  5.740000 2.165000 ;
      RECT  5.640000  0.305000  6.490000 0.475000 ;
      RECT  5.820000  0.895000  6.150000 1.015000 ;
      RECT  5.910000  1.575000  7.850000 1.745000 ;
      RECT  5.920000  2.255000  6.340000 2.635000 ;
      RECT  6.320000  0.475000  6.490000 1.235000 ;
      RECT  6.540000  2.085000  6.780000 2.375000 ;
      RECT  6.670000  0.085000  7.330000 0.565000 ;
      RECT  7.010000  1.945000  7.340000 2.635000 ;
      RECT  7.140000  1.175000  7.470000 1.235000 ;
      RECT  7.510000  0.350000  7.850000 0.680000 ;
      RECT  7.510000  1.745000  7.850000 1.765000 ;
      RECT  7.510000  1.765000  7.680000 2.375000 ;
      RECT  7.640000  0.680000  7.850000 1.575000 ;
      RECT  7.950000  1.915000  8.280000 2.425000 ;
      RECT  8.030000  0.345000  8.280000 1.055000 ;
      RECT  8.030000  1.055000 10.555000 1.275000 ;
      RECT  8.030000  1.275000  8.280000 1.915000 ;
      RECT  8.460000  0.085000  8.745000 0.545000 ;
      RECT  8.460000  1.835000  8.745000 2.635000 ;
      RECT  9.340000  0.085000  9.595000 0.545000 ;
      RECT  9.340000  1.810000  9.595000 2.635000 ;
      RECT 10.105000  0.085000 10.435000 0.545000 ;
      RECT 10.105000  1.810000 10.435000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.615000  1.785000  0.785000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  0.765000  1.235000 0.935000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  1.785000  2.615000 1.955000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  0.765000  3.075000 0.935000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.225000  1.105000  5.395000 1.275000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 0.555000 1.755000 0.845000 1.800000 ;
      RECT 0.555000 1.800000 5.435000 1.940000 ;
      RECT 0.555000 1.940000 0.845000 1.985000 ;
      RECT 1.005000 0.735000 1.295000 0.780000 ;
      RECT 1.005000 0.780000 3.135000 0.920000 ;
      RECT 1.005000 0.920000 1.295000 0.965000 ;
      RECT 2.385000 1.755000 2.675000 1.800000 ;
      RECT 2.385000 1.940000 2.675000 1.985000 ;
      RECT 2.845000 0.735000 3.135000 0.780000 ;
      RECT 2.845000 0.920000 3.135000 0.965000 ;
      RECT 2.920000 0.965000 3.135000 1.120000 ;
      RECT 2.920000 1.120000 5.455000 1.260000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 5.165000 1.075000 5.455000 1.120000 ;
      RECT 5.165000 1.260000 5.455000 1.305000 ;
  END
END sky130_fd_sc_hd__dfstp_4
MACRO sky130_fd_sc_hd__dfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.370000 0.715000 1.650000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.890000 1.495000 7.300000 1.575000 ;
        RECT 6.890000 1.575000 7.220000 2.420000 ;
        RECT 6.900000 0.305000 7.230000 0.740000 ;
        RECT 6.900000 0.740000 7.300000 0.825000 ;
        RECT 7.055000 0.825000 7.300000 0.865000 ;
        RECT 7.065000 1.445000 7.300000 1.495000 ;
        RECT 7.110000 0.865000 7.300000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.315000 1.480000 8.650000 2.465000 ;
        RECT 8.395000 0.255000 8.650000 0.910000 ;
        RECT 8.415000 0.910000 8.650000 1.480000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.930000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.840000 0.805000 ;
      RECT 0.175000  1.795000 0.840000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.200000 2.465000 ;
      RECT 1.440000  2.175000 1.705000 2.635000 ;
      RECT 1.455000  0.085000 1.705000 0.545000 ;
      RECT 1.820000  0.675000 2.045000 0.805000 ;
      RECT 1.820000  0.805000 1.990000 1.910000 ;
      RECT 1.820000  1.910000 2.125000 2.040000 ;
      RECT 1.875000  0.365000 2.210000 0.535000 ;
      RECT 1.875000  0.535000 2.045000 0.675000 ;
      RECT 1.875000  2.040000 2.125000 2.465000 ;
      RECT 2.160000  1.125000 2.400000 1.720000 ;
      RECT 2.215000  0.735000 2.740000 0.955000 ;
      RECT 2.335000  2.190000 3.440000 2.360000 ;
      RECT 2.405000  0.365000 3.080000 0.535000 ;
      RECT 2.570000  0.955000 2.740000 1.655000 ;
      RECT 2.570000  1.655000 3.100000 2.020000 ;
      RECT 2.910000  0.535000 3.080000 1.315000 ;
      RECT 2.910000  1.315000 3.780000 1.485000 ;
      RECT 3.270000  1.485000 3.780000 1.575000 ;
      RECT 3.270000  1.575000 3.440000 2.190000 ;
      RECT 3.290000  0.765000 4.120000 1.065000 ;
      RECT 3.290000  1.065000 3.490000 1.095000 ;
      RECT 3.400000  0.085000 3.770000 0.585000 ;
      RECT 3.610000  1.245000 3.780000 1.315000 ;
      RECT 3.610000  1.835000 3.780000 2.635000 ;
      RECT 3.950000  0.365000 4.355000 0.535000 ;
      RECT 3.950000  0.535000 4.120000 0.765000 ;
      RECT 3.950000  1.065000 4.120000 2.135000 ;
      RECT 3.950000  2.135000 4.200000 2.465000 ;
      RECT 4.290000  1.245000 4.480000 1.965000 ;
      RECT 4.425000  2.165000 5.310000 2.335000 ;
      RECT 4.505000  0.705000 4.970000 1.035000 ;
      RECT 4.525000  0.365000 5.310000 0.535000 ;
      RECT 4.650000  1.035000 4.970000 1.995000 ;
      RECT 5.140000  0.535000 5.310000 0.995000 ;
      RECT 5.140000  0.995000 6.020000 1.325000 ;
      RECT 5.140000  1.325000 5.310000 2.165000 ;
      RECT 5.480000  1.530000 6.380000 1.905000 ;
      RECT 5.490000  2.135000 5.805000 2.635000 ;
      RECT 5.585000  0.085000 5.795000 0.615000 ;
      RECT 6.040000  1.905000 6.380000 2.465000 ;
      RECT 6.060000  0.300000 6.390000 0.825000 ;
      RECT 6.190000  0.825000 6.390000 0.995000 ;
      RECT 6.190000  0.995000 6.940000 1.325000 ;
      RECT 6.190000  1.325000 6.380000 1.530000 ;
      RECT 6.550000  1.625000 6.720000 2.635000 ;
      RECT 6.560000  0.085000 6.730000 0.695000 ;
      RECT 7.410000  1.715000 7.740000 2.445000 ;
      RECT 7.420000  0.345000 7.670000 0.615000 ;
      RECT 7.470000  0.615000 7.670000 0.995000 ;
      RECT 7.470000  0.995000 8.245000 1.325000 ;
      RECT 7.470000  1.325000 7.740000 1.715000 ;
      RECT 7.905000  0.085000 8.225000 0.545000 ;
      RECT 7.930000  1.495000 8.145000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.630000  1.785000 0.800000 1.955000 ;
      RECT 1.025000  1.445000 1.195000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.215000  1.445000 2.385000 1.615000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.730000  1.785000 2.900000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.300000  1.785000 4.470000 1.955000 ;
      RECT 4.735000  1.445000 4.905000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
    LAYER met1 ;
      RECT 0.570000 1.755000 0.860000 1.800000 ;
      RECT 0.570000 1.800000 4.530000 1.940000 ;
      RECT 0.570000 1.940000 0.860000 1.985000 ;
      RECT 0.965000 1.415000 1.255000 1.460000 ;
      RECT 0.965000 1.460000 4.965000 1.600000 ;
      RECT 0.965000 1.600000 1.255000 1.645000 ;
      RECT 2.155000 1.415000 2.445000 1.460000 ;
      RECT 2.155000 1.600000 2.445000 1.645000 ;
      RECT 2.670000 1.755000 2.960000 1.800000 ;
      RECT 2.670000 1.940000 2.960000 1.985000 ;
      RECT 4.240000 1.755000 4.530000 1.800000 ;
      RECT 4.240000 1.940000 4.530000 1.985000 ;
      RECT 4.675000 1.415000 4.965000 1.460000 ;
      RECT 4.675000 1.600000 4.965000 1.645000 ;
  END
END sky130_fd_sc_hd__dfxbp_1
MACRO sky130_fd_sc_hd__dfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.370000 0.715000 1.650000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.890000 1.495000 7.300000 1.575000 ;
        RECT 6.890000 1.575000 7.220000 2.420000 ;
        RECT 6.900000 0.305000 7.230000 0.740000 ;
        RECT 6.900000 0.740000 7.300000 0.825000 ;
        RECT 7.055000 0.825000 7.300000 0.865000 ;
        RECT 7.065000 1.445000 7.300000 1.495000 ;
        RECT 7.110000 0.865000 7.300000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.810000 1.495000 9.145000 2.465000 ;
        RECT 8.890000 0.265000 9.145000 0.885000 ;
        RECT 8.930000 0.885000 9.145000 1.495000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.840000 0.805000 ;
      RECT 0.175000  1.795000 0.840000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.200000 2.465000 ;
      RECT 1.440000  2.175000 1.705000 2.635000 ;
      RECT 1.455000  0.085000 1.705000 0.545000 ;
      RECT 1.820000  0.675000 2.045000 0.805000 ;
      RECT 1.820000  0.805000 1.990000 1.910000 ;
      RECT 1.820000  1.910000 2.125000 2.040000 ;
      RECT 1.875000  0.365000 2.210000 0.535000 ;
      RECT 1.875000  0.535000 2.045000 0.675000 ;
      RECT 1.875000  2.040000 2.125000 2.465000 ;
      RECT 2.160000  1.125000 2.400000 1.720000 ;
      RECT 2.215000  0.735000 2.740000 0.955000 ;
      RECT 2.335000  2.190000 3.440000 2.360000 ;
      RECT 2.405000  0.365000 3.080000 0.535000 ;
      RECT 2.570000  0.955000 2.740000 1.655000 ;
      RECT 2.570000  1.655000 3.100000 2.020000 ;
      RECT 2.910000  0.535000 3.080000 1.315000 ;
      RECT 2.910000  1.315000 3.780000 1.485000 ;
      RECT 3.270000  1.485000 3.780000 1.575000 ;
      RECT 3.270000  1.575000 3.440000 2.190000 ;
      RECT 3.290000  0.765000 4.120000 1.065000 ;
      RECT 3.290000  1.065000 3.490000 1.095000 ;
      RECT 3.400000  0.085000 3.770000 0.585000 ;
      RECT 3.610000  1.245000 3.780000 1.315000 ;
      RECT 3.610000  1.835000 3.780000 2.635000 ;
      RECT 3.950000  0.365000 4.355000 0.535000 ;
      RECT 3.950000  0.535000 4.120000 0.765000 ;
      RECT 3.950000  1.065000 4.120000 2.135000 ;
      RECT 3.950000  2.135000 4.200000 2.465000 ;
      RECT 4.290000  1.245000 4.480000 1.965000 ;
      RECT 4.425000  2.165000 5.310000 2.335000 ;
      RECT 4.505000  0.705000 4.970000 1.035000 ;
      RECT 4.525000  0.365000 5.310000 0.535000 ;
      RECT 4.650000  1.035000 4.970000 1.995000 ;
      RECT 5.140000  0.535000 5.310000 0.995000 ;
      RECT 5.140000  0.995000 6.020000 1.325000 ;
      RECT 5.140000  1.325000 5.310000 2.165000 ;
      RECT 5.480000  1.530000 6.380000 1.905000 ;
      RECT 5.490000  2.135000 5.805000 2.635000 ;
      RECT 5.585000  0.085000 5.795000 0.615000 ;
      RECT 6.040000  1.905000 6.380000 2.465000 ;
      RECT 6.060000  0.300000 6.390000 0.825000 ;
      RECT 6.190000  0.825000 6.390000 0.995000 ;
      RECT 6.190000  0.995000 6.940000 1.325000 ;
      RECT 6.190000  1.325000 6.380000 1.530000 ;
      RECT 6.550000  1.625000 6.720000 2.635000 ;
      RECT 6.560000  0.085000 6.730000 0.695000 ;
      RECT 7.390000  1.720000 7.565000 2.635000 ;
      RECT 7.400000  0.085000 7.570000 0.600000 ;
      RECT 7.905000  0.345000 8.165000 0.615000 ;
      RECT 7.905000  1.715000 8.235000 2.445000 ;
      RECT 7.965000  0.615000 8.165000 0.995000 ;
      RECT 7.965000  0.995000 8.760000 1.325000 ;
      RECT 7.965000  1.325000 8.235000 1.715000 ;
      RECT 8.390000  0.085000 8.720000 0.825000 ;
      RECT 8.425000  1.495000 8.640000 2.635000 ;
      RECT 9.315000  0.085000 9.565000 0.905000 ;
      RECT 9.315000  1.495000 9.565000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.630000  1.785000 0.800000 1.955000 ;
      RECT 1.025000  1.445000 1.195000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.215000  1.445000 2.385000 1.615000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.730000  1.785000 2.900000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.300000  1.785000 4.470000 1.955000 ;
      RECT 4.735000  1.445000 4.905000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 0.570000 1.755000 0.860000 1.800000 ;
      RECT 0.570000 1.800000 4.530000 1.940000 ;
      RECT 0.570000 1.940000 0.860000 1.985000 ;
      RECT 0.965000 1.415000 1.255000 1.460000 ;
      RECT 0.965000 1.460000 4.965000 1.600000 ;
      RECT 0.965000 1.600000 1.255000 1.645000 ;
      RECT 2.155000 1.415000 2.445000 1.460000 ;
      RECT 2.155000 1.600000 2.445000 1.645000 ;
      RECT 2.670000 1.755000 2.960000 1.800000 ;
      RECT 2.670000 1.940000 2.960000 1.985000 ;
      RECT 4.240000 1.755000 4.530000 1.800000 ;
      RECT 4.240000 1.940000 4.530000 1.985000 ;
      RECT 4.675000 1.415000 4.965000 1.460000 ;
      RECT 4.675000 1.600000 4.965000 1.645000 ;
  END
END sky130_fd_sc_hd__dfxbp_2
MACRO sky130_fd_sc_hd__dfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.370000 0.715000 1.650000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.885000 1.495000 7.275000 1.575000 ;
        RECT 6.885000 1.575000 7.215000 2.420000 ;
        RECT 6.895000 0.305000 7.225000 0.740000 ;
        RECT 6.895000 0.740000 7.275000 0.825000 ;
        RECT 7.050000 0.825000 7.275000 0.865000 ;
        RECT 7.060000 1.445000 7.275000 1.495000 ;
        RECT 7.105000 0.865000 7.275000 1.445000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.840000 0.805000 ;
      RECT 0.175000  1.795000 0.840000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.200000 2.465000 ;
      RECT 1.440000  2.175000 1.705000 2.635000 ;
      RECT 1.455000  0.085000 1.705000 0.545000 ;
      RECT 1.820000  0.675000 2.045000 0.805000 ;
      RECT 1.820000  0.805000 1.990000 1.910000 ;
      RECT 1.820000  1.910000 2.125000 2.040000 ;
      RECT 1.875000  0.365000 2.210000 0.535000 ;
      RECT 1.875000  0.535000 2.045000 0.675000 ;
      RECT 1.875000  2.040000 2.125000 2.465000 ;
      RECT 2.160000  1.125000 2.400000 1.720000 ;
      RECT 2.215000  0.735000 2.740000 0.955000 ;
      RECT 2.335000  2.190000 3.440000 2.360000 ;
      RECT 2.405000  0.365000 3.080000 0.535000 ;
      RECT 2.570000  0.955000 2.740000 1.655000 ;
      RECT 2.570000  1.655000 3.100000 2.020000 ;
      RECT 2.910000  0.535000 3.080000 1.315000 ;
      RECT 2.910000  1.315000 3.780000 1.485000 ;
      RECT 3.270000  1.485000 3.780000 1.575000 ;
      RECT 3.270000  1.575000 3.440000 2.190000 ;
      RECT 3.290000  0.765000 4.120000 1.065000 ;
      RECT 3.290000  1.065000 3.490000 1.095000 ;
      RECT 3.400000  0.085000 3.770000 0.585000 ;
      RECT 3.610000  1.245000 3.780000 1.315000 ;
      RECT 3.610000  1.835000 3.780000 2.635000 ;
      RECT 3.950000  0.365000 4.355000 0.535000 ;
      RECT 3.950000  0.535000 4.120000 0.765000 ;
      RECT 3.950000  1.065000 4.120000 2.135000 ;
      RECT 3.950000  2.135000 4.200000 2.465000 ;
      RECT 4.290000  1.245000 4.480000 1.965000 ;
      RECT 4.425000  2.165000 5.310000 2.335000 ;
      RECT 4.505000  0.705000 4.970000 1.035000 ;
      RECT 4.525000  0.365000 5.310000 0.535000 ;
      RECT 4.650000  1.035000 4.970000 1.995000 ;
      RECT 5.140000  0.535000 5.310000 0.995000 ;
      RECT 5.140000  0.995000 6.015000 1.325000 ;
      RECT 5.140000  1.325000 5.310000 2.165000 ;
      RECT 5.480000  1.530000 6.375000 1.905000 ;
      RECT 5.490000  2.135000 5.805000 2.635000 ;
      RECT 5.585000  0.085000 5.795000 0.615000 ;
      RECT 6.035000  1.905000 6.375000 2.465000 ;
      RECT 6.055000  0.300000 6.385000 0.825000 ;
      RECT 6.185000  0.825000 6.385000 0.995000 ;
      RECT 6.185000  0.995000 6.935000 1.325000 ;
      RECT 6.185000  1.325000 6.375000 1.530000 ;
      RECT 6.545000  1.625000 6.715000 2.635000 ;
      RECT 6.555000  0.085000 6.725000 0.695000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.630000  1.785000 0.800000 1.955000 ;
      RECT 1.025000  1.445000 1.195000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.215000  1.445000 2.385000 1.615000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.730000  1.785000 2.900000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.300000  1.785000 4.470000 1.955000 ;
      RECT 4.735000  1.445000 4.905000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
    LAYER met1 ;
      RECT 0.570000 1.755000 0.860000 1.800000 ;
      RECT 0.570000 1.800000 4.530000 1.940000 ;
      RECT 0.570000 1.940000 0.860000 1.985000 ;
      RECT 0.965000 1.415000 1.255000 1.460000 ;
      RECT 0.965000 1.460000 4.965000 1.600000 ;
      RECT 0.965000 1.600000 1.255000 1.645000 ;
      RECT 2.155000 1.415000 2.445000 1.460000 ;
      RECT 2.155000 1.600000 2.445000 1.645000 ;
      RECT 2.670000 1.755000 2.960000 1.800000 ;
      RECT 2.670000 1.940000 2.960000 1.985000 ;
      RECT 4.240000 1.755000 4.530000 1.800000 ;
      RECT 4.240000 1.940000 4.530000 1.985000 ;
      RECT 4.675000 1.415000 4.965000 1.460000 ;
      RECT 4.675000 1.600000 4.965000 1.645000 ;
  END
END sky130_fd_sc_hd__dfxtp_1
MACRO sky130_fd_sc_hd__dfxtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.370000 0.715000 1.650000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.885000 1.495000 7.275000 1.575000 ;
        RECT 6.885000 1.575000 7.215000 2.420000 ;
        RECT 6.895000 0.305000 7.225000 0.740000 ;
        RECT 6.895000 0.740000 7.275000 0.825000 ;
        RECT 7.050000 0.825000 7.275000 0.865000 ;
        RECT 7.060000 1.445000 7.275000 1.495000 ;
        RECT 7.105000 0.865000 7.275000 1.445000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.840000 0.805000 ;
      RECT 0.175000  1.795000 0.840000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.200000 2.465000 ;
      RECT 1.440000  2.175000 1.705000 2.635000 ;
      RECT 1.455000  0.085000 1.705000 0.545000 ;
      RECT 1.820000  0.675000 2.045000 0.805000 ;
      RECT 1.820000  0.805000 1.990000 1.910000 ;
      RECT 1.820000  1.910000 2.125000 2.040000 ;
      RECT 1.875000  0.365000 2.210000 0.535000 ;
      RECT 1.875000  0.535000 2.045000 0.675000 ;
      RECT 1.875000  2.040000 2.125000 2.465000 ;
      RECT 2.160000  1.125000 2.400000 1.720000 ;
      RECT 2.215000  0.735000 2.740000 0.955000 ;
      RECT 2.335000  2.190000 3.440000 2.360000 ;
      RECT 2.405000  0.365000 3.080000 0.535000 ;
      RECT 2.570000  0.955000 2.740000 1.655000 ;
      RECT 2.570000  1.655000 3.100000 2.020000 ;
      RECT 2.910000  0.535000 3.080000 1.315000 ;
      RECT 2.910000  1.315000 3.780000 1.485000 ;
      RECT 3.270000  1.485000 3.780000 1.575000 ;
      RECT 3.270000  1.575000 3.440000 2.190000 ;
      RECT 3.290000  0.765000 4.120000 1.065000 ;
      RECT 3.290000  1.065000 3.490000 1.095000 ;
      RECT 3.400000  0.085000 3.770000 0.585000 ;
      RECT 3.610000  1.245000 3.780000 1.315000 ;
      RECT 3.610000  1.835000 3.780000 2.635000 ;
      RECT 3.950000  0.365000 4.355000 0.535000 ;
      RECT 3.950000  0.535000 4.120000 0.765000 ;
      RECT 3.950000  1.065000 4.120000 2.135000 ;
      RECT 3.950000  2.135000 4.200000 2.465000 ;
      RECT 4.290000  1.245000 4.480000 1.965000 ;
      RECT 4.425000  2.165000 5.310000 2.335000 ;
      RECT 4.505000  0.705000 4.970000 1.035000 ;
      RECT 4.525000  0.365000 5.310000 0.535000 ;
      RECT 4.650000  1.035000 4.970000 1.995000 ;
      RECT 5.140000  0.535000 5.310000 0.995000 ;
      RECT 5.140000  0.995000 6.015000 1.325000 ;
      RECT 5.140000  1.325000 5.310000 2.165000 ;
      RECT 5.480000  1.530000 6.375000 1.905000 ;
      RECT 5.490000  2.135000 5.805000 2.635000 ;
      RECT 5.585000  0.085000 5.795000 0.615000 ;
      RECT 6.035000  1.905000 6.375000 2.465000 ;
      RECT 6.055000  0.300000 6.385000 0.825000 ;
      RECT 6.185000  0.825000 6.385000 0.995000 ;
      RECT 6.185000  0.995000 6.935000 1.325000 ;
      RECT 6.185000  1.325000 6.375000 1.530000 ;
      RECT 6.545000  1.625000 6.715000 2.635000 ;
      RECT 6.555000  0.085000 6.725000 0.695000 ;
      RECT 7.385000  1.720000 7.555000 2.635000 ;
      RECT 7.395000  0.085000 7.565000 0.600000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.630000  1.785000 0.800000 1.955000 ;
      RECT 1.025000  1.445000 1.195000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.215000  1.445000 2.385000 1.615000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.730000  1.785000 2.900000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.300000  1.785000 4.470000 1.955000 ;
      RECT 4.735000  1.445000 4.905000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 0.570000 1.755000 0.860000 1.800000 ;
      RECT 0.570000 1.800000 4.530000 1.940000 ;
      RECT 0.570000 1.940000 0.860000 1.985000 ;
      RECT 0.965000 1.415000 1.255000 1.460000 ;
      RECT 0.965000 1.460000 4.965000 1.600000 ;
      RECT 0.965000 1.600000 1.255000 1.645000 ;
      RECT 2.155000 1.415000 2.445000 1.460000 ;
      RECT 2.155000 1.600000 2.445000 1.645000 ;
      RECT 2.670000 1.755000 2.960000 1.800000 ;
      RECT 2.670000 1.940000 2.960000 1.985000 ;
      RECT 4.240000 1.755000 4.530000 1.800000 ;
      RECT 4.240000 1.940000 4.530000 1.985000 ;
      RECT 4.675000 1.415000 4.965000 1.460000 ;
      RECT 4.675000 1.600000 4.965000 1.645000 ;
  END
END sky130_fd_sc_hd__dfxtp_2
MACRO sky130_fd_sc_hd__dfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.440000 1.065000 1.720000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.985000 0.305000 7.320000 0.730000 ;
        RECT 6.985000 0.730000 8.655000 0.900000 ;
        RECT 6.985000 1.465000 8.655000 1.635000 ;
        RECT 6.985000 1.635000 7.320000 2.395000 ;
        RECT 7.840000 0.305000 8.175000 0.730000 ;
        RECT 7.840000 1.635000 8.170000 2.395000 ;
        RECT 8.410000 0.900000 8.655000 1.465000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.930000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.840000 0.805000 ;
      RECT 0.175000  1.795000 0.840000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.240000 2.465000 ;
      RECT 1.440000  2.175000 1.705000 2.635000 ;
      RECT 1.455000  0.085000 1.705000 0.545000 ;
      RECT 1.890000  0.365000 2.220000 0.535000 ;
      RECT 1.890000  0.535000 2.060000 2.065000 ;
      RECT 1.890000  2.065000 2.125000 2.440000 ;
      RECT 2.230000  0.705000 2.810000 1.035000 ;
      RECT 2.230000  1.035000 2.470000 1.905000 ;
      RECT 2.370000  2.190000 3.440000 2.360000 ;
      RECT 2.400000  0.365000 3.150000 0.535000 ;
      RECT 2.660000  1.655000 3.100000 2.010000 ;
      RECT 2.980000  0.535000 3.150000 1.315000 ;
      RECT 2.980000  1.315000 3.780000 1.485000 ;
      RECT 3.270000  1.485000 3.780000 1.575000 ;
      RECT 3.270000  1.575000 3.440000 2.190000 ;
      RECT 3.320000  0.765000 4.120000 1.065000 ;
      RECT 3.320000  1.065000 3.490000 1.095000 ;
      RECT 3.400000  0.085000 3.770000 0.585000 ;
      RECT 3.610000  1.245000 3.780000 1.315000 ;
      RECT 3.610000  1.835000 3.780000 2.635000 ;
      RECT 3.950000  0.365000 4.410000 0.535000 ;
      RECT 3.950000  0.535000 4.120000 0.765000 ;
      RECT 3.950000  1.065000 4.120000 2.135000 ;
      RECT 3.950000  2.135000 4.200000 2.465000 ;
      RECT 4.290000  0.705000 4.840000 1.035000 ;
      RECT 4.290000  1.245000 4.480000 1.965000 ;
      RECT 4.425000  2.165000 5.310000 2.335000 ;
      RECT 4.640000  0.365000 5.310000 0.535000 ;
      RECT 4.650000  1.035000 4.840000 1.575000 ;
      RECT 4.650000  1.575000 4.970000 1.905000 ;
      RECT 5.140000  0.535000 5.310000 1.075000 ;
      RECT 5.140000  1.075000 6.230000 1.245000 ;
      RECT 5.140000  1.245000 5.310000 2.165000 ;
      RECT 5.480000  1.500000 6.590000 1.670000 ;
      RECT 5.480000  1.670000 6.340000 1.830000 ;
      RECT 5.490000  2.135000 5.705000 2.635000 ;
      RECT 5.625000  0.085000 5.795000 0.615000 ;
      RECT 6.090000  0.295000 6.450000 0.735000 ;
      RECT 6.090000  0.735000 6.590000 0.905000 ;
      RECT 6.170000  1.830000 6.340000 2.455000 ;
      RECT 6.420000  0.905000 6.590000 1.075000 ;
      RECT 6.420000  1.075000 8.240000 1.245000 ;
      RECT 6.420000  1.245000 6.590000 1.500000 ;
      RECT 6.625000  0.085000 6.795000 0.565000 ;
      RECT 6.625000  1.855000 6.805000 2.635000 ;
      RECT 7.495000  0.085000 7.665000 0.560000 ;
      RECT 7.500000  1.805000 7.670000 2.635000 ;
      RECT 8.340000  1.805000 8.510000 2.635000 ;
      RECT 8.345000  0.085000 8.515000 0.560000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.785000 0.780000 1.955000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  0.765000 1.240000 0.935000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  0.765000 2.640000 0.935000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  1.785000 3.100000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.310000  0.765000 4.480000 0.935000 ;
      RECT 4.310000  1.785000 4.480000 1.955000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.755000 0.840000 1.800000 ;
      RECT 0.550000 1.800000 4.540000 1.940000 ;
      RECT 0.550000 1.940000 0.840000 1.985000 ;
      RECT 1.010000 0.735000 1.300000 0.780000 ;
      RECT 1.010000 0.780000 4.540000 0.920000 ;
      RECT 1.010000 0.920000 1.300000 0.965000 ;
      RECT 2.410000 0.735000 2.700000 0.780000 ;
      RECT 2.410000 0.920000 2.700000 0.965000 ;
      RECT 2.870000 1.755000 3.160000 1.800000 ;
      RECT 2.870000 1.940000 3.160000 1.985000 ;
      RECT 4.250000 0.735000 4.540000 0.780000 ;
      RECT 4.250000 0.920000 4.540000 0.965000 ;
      RECT 4.250000 1.755000 4.540000 1.800000 ;
      RECT 4.250000 1.940000 4.540000 1.985000 ;
  END
END sky130_fd_sc_hd__dfxtp_4
MACRO sky130_fd_sc_hd__diode_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__diode_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.920000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DIODE
    ANTENNADIFFAREA  0.434700 ;
    ANTENNAGATEAREA  0.434700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.835000 2.465000 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.920000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.110000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.920000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.920000 0.085000 ;
      RECT 0.000000  2.635000 0.920000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
  END
END sky130_fd_sc_hd__diode_2
MACRO sky130_fd_sc_hd__dlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlclkp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 1.435000 2.185000 1.685000 ;
        RECT 1.985000 0.385000 2.185000 1.435000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.055000 0.255000 6.355000 0.595000 ;
        RECT 6.090000 1.495000 6.355000 2.455000 ;
        RECT 6.170000 0.595000 6.355000 1.495000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
      LAYER mcon ;
        RECT 0.145000 1.105000 0.315000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.190000 1.105000 5.510000 1.435000 ;
      LAYER mcon ;
        RECT 5.210000 1.105000 5.380000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.085000 1.075000 0.380000 1.120000 ;
        RECT 0.085000 1.120000 5.440000 1.260000 ;
        RECT 0.085000 1.260000 0.380000 1.305000 ;
        RECT 5.150000 1.075000 5.440000 1.120000 ;
        RECT 5.150000 1.260000 5.440000 1.305000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 0.995000 1.355000 ;
        RECT -0.190000 1.355000 6.630000 2.910000 ;
        RECT  2.620000 1.305000 6.630000 1.355000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.175000  0.260000 0.345000 0.615000 ;
      RECT 0.175000  0.615000 0.780000 0.785000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.445000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.785000 0.780000 1.060000 ;
      RECT 0.610000  1.060000 0.840000 1.390000 ;
      RECT 0.610000  1.390000 0.780000 1.795000 ;
      RECT 1.015000  0.260000 1.280000 1.855000 ;
      RECT 1.015000  1.855000 2.590000 2.025000 ;
      RECT 1.015000  2.025000 1.240000 2.465000 ;
      RECT 1.450000  2.195000 1.815000 2.635000 ;
      RECT 1.480000  0.085000 1.810000 0.905000 ;
      RECT 2.390000  0.815000 3.220000 0.985000 ;
      RECT 2.390000  0.985000 2.590000 1.855000 ;
      RECT 2.475000  2.255000 3.225000 2.425000 ;
      RECT 2.790000  0.390000 3.725000 0.560000 ;
      RECT 3.055000  1.155000 4.175000 1.325000 ;
      RECT 3.055000  1.325000 3.225000 2.255000 ;
      RECT 3.395000  2.135000 3.695000 2.635000 ;
      RECT 3.430000  1.535000 4.710000 1.840000 ;
      RECT 3.430000  1.840000 4.130000 1.865000 ;
      RECT 3.555000  0.560000 3.725000 0.995000 ;
      RECT 3.555000  0.995000 4.175000 1.155000 ;
      RECT 3.895000  0.085000 4.145000 0.610000 ;
      RECT 3.910000  1.865000 4.130000 2.435000 ;
      RECT 4.310000  2.010000 4.595000 2.635000 ;
      RECT 4.320000  0.255000 4.580000 0.615000 ;
      RECT 4.345000  0.615000 4.580000 0.995000 ;
      RECT 4.345000  0.995000 4.740000 1.325000 ;
      RECT 4.345000  1.325000 4.710000 1.535000 ;
      RECT 4.840000  0.290000 5.155000 0.620000 ;
      RECT 4.935000  0.620000 5.155000 0.765000 ;
      RECT 4.935000  0.765000 6.000000 0.935000 ;
      RECT 5.005000  1.725000 5.920000 1.895000 ;
      RECT 5.005000  1.895000 5.335000 2.465000 ;
      RECT 5.570000  2.130000 5.920000 2.635000 ;
      RECT 5.670000  0.085000 5.840000 0.545000 ;
      RECT 5.750000  0.935000 6.000000 1.325000 ;
      RECT 5.750000  1.325000 5.920000 1.725000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__dlclkp_1
MACRO sky130_fd_sc_hd__dlclkp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlclkp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 1.435000 2.215000 1.685000 ;
        RECT 1.985000 0.285000 2.215000 1.435000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.060000 0.255000 6.360000 0.595000 ;
        RECT 6.095000 1.495000 6.360000 2.455000 ;
        RECT 6.165000 0.595000 6.360000 1.495000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.985000 0.330000 1.625000 ;
      LAYER mcon ;
        RECT 0.150000 1.105000 0.320000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.210000 1.105000 5.485000 1.435000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.090000 1.075000 0.380000 1.120000 ;
        RECT 0.090000 1.120000 5.440000 1.260000 ;
        RECT 0.090000 1.260000 0.380000 1.305000 ;
        RECT 5.150000 1.075000 5.440000 1.120000 ;
        RECT 5.150000 1.260000 5.440000 1.305000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 0.995000 1.355000 ;
        RECT -0.190000 1.355000 7.090000 2.910000 ;
        RECT  2.625000 1.305000 7.090000 1.355000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.175000  0.260000 0.345000 0.615000 ;
      RECT 0.175000  0.615000 0.780000 0.785000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.445000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.785000 0.780000 1.060000 ;
      RECT 0.610000  1.060000 0.840000 1.390000 ;
      RECT 0.610000  1.390000 0.780000 1.795000 ;
      RECT 1.015000  0.260000 1.280000 1.855000 ;
      RECT 1.015000  1.855000 2.645000 2.025000 ;
      RECT 1.015000  2.025000 1.240000 2.465000 ;
      RECT 1.455000  2.195000 1.820000 2.635000 ;
      RECT 1.485000  0.085000 1.815000 0.905000 ;
      RECT 2.395000  0.815000 3.225000 0.985000 ;
      RECT 2.395000  0.985000 2.645000 1.855000 ;
      RECT 2.480000  2.255000 3.230000 2.425000 ;
      RECT 2.795000  0.390000 3.725000 0.560000 ;
      RECT 3.060000  1.155000 4.180000 1.325000 ;
      RECT 3.060000  1.325000 3.230000 2.255000 ;
      RECT 3.400000  2.135000 3.700000 2.635000 ;
      RECT 3.435000  1.535000 4.735000 1.840000 ;
      RECT 3.435000  1.840000 4.135000 1.865000 ;
      RECT 3.555000  0.560000 3.725000 0.995000 ;
      RECT 3.555000  0.995000 4.180000 1.155000 ;
      RECT 3.895000  0.085000 4.145000 0.610000 ;
      RECT 3.915000  1.865000 4.135000 2.435000 ;
      RECT 4.315000  0.255000 4.585000 0.615000 ;
      RECT 4.315000  2.010000 4.600000 2.635000 ;
      RECT 4.350000  0.615000 4.585000 0.995000 ;
      RECT 4.350000  0.995000 4.735000 1.535000 ;
      RECT 4.835000  0.290000 5.150000 0.620000 ;
      RECT 4.930000  0.620000 5.150000 0.765000 ;
      RECT 4.930000  0.765000 5.995000 0.935000 ;
      RECT 5.010000  1.725000 5.925000 1.895000 ;
      RECT 5.010000  1.895000 5.340000 2.465000 ;
      RECT 5.575000  2.130000 5.925000 2.635000 ;
      RECT 5.675000  0.085000 5.845000 0.545000 ;
      RECT 5.755000  0.935000 5.995000 1.325000 ;
      RECT 5.755000  1.325000 5.925000 1.725000 ;
      RECT 6.530000  0.085000 6.810000 0.885000 ;
      RECT 6.530000  1.485000 6.810000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
END sky130_fd_sc_hd__dlclkp_2
MACRO sky130_fd_sc_hd__dlclkp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlclkp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 0.765000 1.950000 1.015000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  1.039500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.040000 0.255000 6.460000 0.545000 ;
        RECT 6.040000 1.835000 7.300000 2.005000 ;
        RECT 6.040000 2.005000 6.370000 2.455000 ;
        RECT 6.290000 0.545000 6.460000 0.715000 ;
        RECT 6.290000 0.715000 7.300000 0.885000 ;
        RECT 6.585000 1.785000 7.300000 1.835000 ;
        RECT 6.750000 0.885000 7.300000 1.785000 ;
        RECT 6.970000 0.255000 7.300000 0.715000 ;
        RECT 6.970000 2.005000 7.300000 2.465000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.406500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.985000 0.330000 1.625000 ;
      LAYER mcon ;
        RECT 0.150000 1.105000 0.320000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.230000 1.055000 5.740000 1.325000 ;
      LAYER mcon ;
        RECT 5.230000 1.105000 5.400000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.090000 1.075000 0.380000 1.120000 ;
        RECT 0.090000 1.120000 5.460000 1.260000 ;
        RECT 0.090000 1.260000 0.380000 1.305000 ;
        RECT 5.170000 1.075000 5.460000 1.120000 ;
        RECT 5.170000 1.260000 5.460000 1.305000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.635000 ;
      RECT 0.085000  0.635000 0.780000 0.805000 ;
      RECT 0.085000  1.795000 0.780000 1.965000 ;
      RECT 0.085000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.280000 1.355000 ;
      RECT 1.015000  1.355000 2.335000 1.585000 ;
      RECT 1.015000  1.585000 1.240000 2.465000 ;
      RECT 1.450000  0.085000 1.785000 0.465000 ;
      RECT 1.450000  2.195000 1.815000 2.635000 ;
      RECT 1.525000  1.785000 1.695000 1.855000 ;
      RECT 1.525000  1.855000 2.845000 1.905000 ;
      RECT 1.525000  1.905000 2.735000 2.025000 ;
      RECT 2.045000  1.585000 2.335000 1.685000 ;
      RECT 2.290000  0.705000 2.735000 1.035000 ;
      RECT 2.415000  0.365000 3.075000 0.535000 ;
      RECT 2.475000  2.195000 3.165000 2.425000 ;
      RECT 2.505000  1.575000 2.845000 1.855000 ;
      RECT 2.565000  1.035000 2.735000 1.575000 ;
      RECT 2.905000  0.535000 3.075000 0.995000 ;
      RECT 2.905000  0.995000 3.775000 1.165000 ;
      RECT 2.915000  2.060000 3.185000 2.090000 ;
      RECT 2.915000  2.090000 3.180000 2.105000 ;
      RECT 2.915000  2.105000 3.165000 2.195000 ;
      RECT 2.980000  2.015000 3.185000 2.060000 ;
      RECT 3.015000  1.165000 3.775000 1.325000 ;
      RECT 3.015000  1.325000 3.185000 2.015000 ;
      RECT 3.315000  0.085000 3.650000 0.530000 ;
      RECT 3.335000  2.175000 3.695000 2.635000 ;
      RECT 3.355000  1.535000 4.115000 1.865000 ;
      RECT 3.895000  0.415000 4.115000 0.745000 ;
      RECT 3.895000  1.865000 4.115000 2.435000 ;
      RECT 3.945000  0.745000 4.115000 0.995000 ;
      RECT 3.945000  0.995000 4.720000 1.325000 ;
      RECT 3.945000  1.325000 4.115000 1.535000 ;
      RECT 4.295000  0.085000 4.580000 0.715000 ;
      RECT 4.295000  2.010000 4.580000 2.635000 ;
      RECT 4.750000  0.290000 5.060000 0.715000 ;
      RECT 4.750000  0.715000 6.120000 0.825000 ;
      RECT 4.750000  1.495000 6.140000 1.665000 ;
      RECT 4.750000  1.665000 5.035000 2.465000 ;
      RECT 4.890000  0.825000 6.120000 0.885000 ;
      RECT 4.890000  0.885000 5.060000 1.495000 ;
      RECT 5.575000  1.835000 5.840000 2.635000 ;
      RECT 5.590000  0.085000 5.870000 0.545000 ;
      RECT 5.910000  0.885000 6.120000 1.055000 ;
      RECT 5.910000  1.055000 6.580000 1.290000 ;
      RECT 5.910000  1.290000 6.140000 1.495000 ;
      RECT 6.540000  2.175000 6.800000 2.635000 ;
      RECT 6.630000  0.085000 6.800000 0.545000 ;
      RECT 7.470000  0.085000 7.735000 0.885000 ;
      RECT 7.470000  1.485000 7.735000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.785000 0.780000 1.955000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.755000 0.840000 1.800000 ;
      RECT 0.550000 1.800000 1.755000 1.940000 ;
      RECT 0.550000 1.940000 0.840000 1.985000 ;
      RECT 1.465000 1.755000 1.755000 1.800000 ;
      RECT 1.465000 1.940000 1.755000 1.985000 ;
  END
END sky130_fd_sc_hd__dlclkp_4
MACRO sky130_fd_sc_hd__dlrbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.060000 0.255000 6.380000 2.465000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.475000 0.255000 7.735000 0.595000 ;
        RECT 7.475000 1.785000 7.735000 2.465000 ;
        RECT 7.560000 0.595000 7.735000 1.785000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.470000 0.995000 5.455000 1.325000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.635000 ;
      RECT 0.085000  0.635000 0.780000 0.805000 ;
      RECT 0.085000  1.795000 0.780000 1.965000 ;
      RECT 0.085000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.455000  1.495000 2.140000 1.665000 ;
      RECT 1.455000  1.665000 1.785000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.140000 0.765000 ;
      RECT 1.535000  0.765000 2.340000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.955000  1.835000 2.270000 2.635000 ;
      RECT 1.970000  0.785000 2.340000 1.095000 ;
      RECT 1.970000  1.095000 2.140000 1.495000 ;
      RECT 2.470000  1.355000 2.755000 2.005000 ;
      RECT 2.715000  0.705000 3.095000 1.035000 ;
      RECT 2.840000  0.365000 3.500000 0.535000 ;
      RECT 2.900000  2.255000 3.650000 2.425000 ;
      RECT 2.925000  1.035000 3.095000 1.415000 ;
      RECT 2.925000  1.415000 3.265000 1.995000 ;
      RECT 3.330000  0.535000 3.500000 0.995000 ;
      RECT 3.330000  0.995000 4.300000 1.165000 ;
      RECT 3.480000  1.165000 4.300000 1.325000 ;
      RECT 3.480000  1.325000 3.650000 2.255000 ;
      RECT 3.740000  0.085000 4.070000 0.530000 ;
      RECT 3.820000  2.135000 4.090000 2.635000 ;
      RECT 3.840000  1.535000 5.875000 1.765000 ;
      RECT 3.840000  1.765000 4.970000 1.865000 ;
      RECT 4.240000  0.255000 4.540000 0.655000 ;
      RECT 4.240000  0.655000 5.875000 0.825000 ;
      RECT 4.260000  2.135000 4.590000 2.635000 ;
      RECT 4.760000  1.865000 4.970000 2.435000 ;
      RECT 5.135000  0.085000 5.875000 0.485000 ;
      RECT 5.150000  1.935000 5.890000 2.635000 ;
      RECT 5.625000  0.825000 5.875000 1.535000 ;
      RECT 6.580000  0.255000 6.750000 0.985000 ;
      RECT 6.580000  0.985000 6.830000 0.995000 ;
      RECT 6.580000  0.995000 7.390000 1.325000 ;
      RECT 6.580000  1.325000 6.830000 2.465000 ;
      RECT 6.975000  0.085000 7.305000 0.465000 ;
      RECT 7.010000  1.835000 7.305000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.785000 2.640000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  1.445000 3.100000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.160000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.700000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.755000 2.700000 1.800000 ;
      RECT 2.410000 1.940000 2.700000 1.985000 ;
      RECT 2.870000 1.415000 3.160000 1.460000 ;
      RECT 2.870000 1.600000 3.160000 1.645000 ;
  END
END sky130_fd_sc_hd__dlrbn_1
MACRO sky130_fd_sc_hd__dlrbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrbn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.536250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.650000 0.415000 5.910000 0.655000 ;
        RECT 5.650000 0.655000 5.950000 0.685000 ;
        RECT 5.650000 0.685000 5.975000 0.825000 ;
        RECT 5.650000 1.495000 5.975000 1.660000 ;
        RECT 5.650000 1.660000 5.915000 2.465000 ;
        RECT 5.740000 0.825000 5.975000 0.860000 ;
        RECT 5.790000 0.860000 5.975000 0.885000 ;
        RECT 5.790000 0.885000 6.355000 1.325000 ;
        RECT 5.790000 1.325000 5.975000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.500000 0.255000 7.755000 0.825000 ;
        RECT 7.500000 1.445000 7.755000 2.465000 ;
        RECT 7.545000 0.825000 7.755000 1.055000 ;
        RECT 7.545000 1.055000 8.195000 1.325000 ;
        RECT 7.545000 1.325000 7.755000 1.445000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.390000 0.995000 5.140000 1.325000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.635000 ;
      RECT 0.085000  0.635000 0.780000 0.805000 ;
      RECT 0.085000  1.795000 0.780000 1.965000 ;
      RECT 0.085000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.605000  0.805000 0.780000 1.070000 ;
      RECT 0.605000  1.070000 0.840000 1.400000 ;
      RECT 0.605000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.455000  1.495000 2.140000 1.665000 ;
      RECT 1.455000  1.665000 1.785000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.140000 0.765000 ;
      RECT 1.535000  0.765000 2.340000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.955000  1.835000 2.270000 2.635000 ;
      RECT 1.970000  0.785000 2.340000 1.095000 ;
      RECT 1.970000  1.095000 2.140000 1.495000 ;
      RECT 2.470000  1.355000 2.755000 2.005000 ;
      RECT 2.715000  0.705000 3.095000 1.035000 ;
      RECT 2.840000  0.365000 3.500000 0.535000 ;
      RECT 2.900000  2.255000 3.650000 2.425000 ;
      RECT 2.925000  1.035000 3.095000 1.415000 ;
      RECT 2.925000  1.415000 3.265000 1.995000 ;
      RECT 3.330000  0.535000 3.500000 0.995000 ;
      RECT 3.330000  0.995000 4.200000 1.165000 ;
      RECT 3.480000  1.165000 4.200000 1.325000 ;
      RECT 3.480000  1.325000 3.650000 2.255000 ;
      RECT 3.740000  0.085000 4.070000 0.825000 ;
      RECT 3.820000  2.135000 4.590000 2.635000 ;
      RECT 3.840000  1.495000 5.480000 1.665000 ;
      RECT 3.840000  1.665000 4.930000 1.865000 ;
      RECT 4.340000  0.415000 4.560000 0.655000 ;
      RECT 4.340000  0.655000 5.480000 0.825000 ;
      RECT 4.760000  1.865000 4.930000 2.435000 ;
      RECT 5.100000  0.085000 5.480000 0.485000 ;
      RECT 5.100000  1.855000 5.350000 2.635000 ;
      RECT 5.310000  0.825000 5.480000 0.995000 ;
      RECT 5.310000  0.995000 5.620000 1.325000 ;
      RECT 5.310000  1.325000 5.480000 1.495000 ;
      RECT 6.085000  0.085000 6.355000 0.545000 ;
      RECT 6.085000  1.830000 6.355000 2.635000 ;
      RECT 6.525000  0.255000 6.855000 0.995000 ;
      RECT 6.525000  0.995000 7.375000 1.325000 ;
      RECT 6.525000  1.325000 6.855000 2.465000 ;
      RECT 7.025000  0.085000 7.330000 0.545000 ;
      RECT 7.035000  1.835000 7.330000 2.635000 ;
      RECT 7.925000  0.085000 8.195000 0.885000 ;
      RECT 7.925000  1.495000 8.195000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.785000 2.640000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  1.445000 3.100000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.160000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.700000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.755000 2.700000 1.800000 ;
      RECT 2.410000 1.940000 2.700000 1.985000 ;
      RECT 2.870000 1.415000 3.160000 1.460000 ;
      RECT 2.870000 1.600000 3.160000 1.645000 ;
  END
END sky130_fd_sc_hd__dlrbn_2
MACRO sky130_fd_sc_hd__dlrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.060000 0.255000 6.410000 2.465000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.475000 0.255000 7.735000 0.595000 ;
        RECT 7.475000 1.785000 7.735000 2.465000 ;
        RECT 7.565000 0.595000 7.735000 1.785000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.450000 0.995000 5.435000 1.325000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.325000 1.625000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.635000 ;
      RECT 0.085000  0.635000 0.780000 0.805000 ;
      RECT 0.085000  1.795000 0.780000 1.965000 ;
      RECT 0.085000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.455000  1.495000 2.140000 1.665000 ;
      RECT 1.455000  1.665000 1.785000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.140000 0.765000 ;
      RECT 1.535000  0.765000 2.340000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.955000  1.835000 2.270000 2.635000 ;
      RECT 1.970000  0.785000 2.340000 1.095000 ;
      RECT 1.970000  1.095000 2.140000 1.495000 ;
      RECT 2.470000  1.355000 2.755000 1.685000 ;
      RECT 2.600000  0.765000 3.095000 1.035000 ;
      RECT 2.745000  2.255000 3.585000 2.425000 ;
      RECT 2.770000  0.365000 3.500000 0.535000 ;
      RECT 2.925000  1.035000 3.095000 1.575000 ;
      RECT 2.925000  1.575000 3.265000 1.905000 ;
      RECT 2.925000  1.905000 3.130000 1.995000 ;
      RECT 3.270000  2.125000 3.585000 2.255000 ;
      RECT 3.305000  2.075000 3.585000 2.125000 ;
      RECT 3.330000  0.535000 3.500000 0.995000 ;
      RECT 3.330000  0.995000 4.200000 1.165000 ;
      RECT 3.395000  2.015000 3.605000 2.045000 ;
      RECT 3.395000  2.045000 3.585000 2.075000 ;
      RECT 3.415000  1.990000 3.605000 2.015000 ;
      RECT 3.420000  1.975000 3.605000 1.990000 ;
      RECT 3.430000  1.960000 3.605000 1.975000 ;
      RECT 3.435000  1.165000 4.200000 1.325000 ;
      RECT 3.435000  1.325000 3.605000 1.960000 ;
      RECT 3.735000  0.085000 4.070000 0.530000 ;
      RECT 3.755000  2.135000 4.590000 2.635000 ;
      RECT 3.840000  1.535000 5.890000 1.765000 ;
      RECT 3.840000  1.765000 4.950000 1.865000 ;
      RECT 4.240000  0.255000 4.540000 0.655000 ;
      RECT 4.240000  0.655000 5.890000 0.825000 ;
      RECT 4.780000  1.865000 4.950000 2.435000 ;
      RECT 5.120000  0.085000 5.890000 0.485000 ;
      RECT 5.120000  1.935000 5.890000 2.635000 ;
      RECT 5.655000  0.825000 5.890000 1.535000 ;
      RECT 6.580000  0.255000 6.805000 0.995000 ;
      RECT 6.580000  0.995000 7.395000 1.325000 ;
      RECT 6.580000  1.325000 6.830000 2.465000 ;
      RECT 6.975000  0.085000 7.305000 0.465000 ;
      RECT 7.010000  1.835000 7.305000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.445000 2.640000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.925000  1.785000 3.095000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 2.700000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 3.155000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.415000 2.700000 1.460000 ;
      RECT 2.410000 1.600000 2.700000 1.645000 ;
      RECT 2.865000 1.755000 3.155000 1.800000 ;
      RECT 2.865000 1.940000 3.155000 1.985000 ;
  END
END sky130_fd_sc_hd__dlrbp_1
MACRO sky130_fd_sc_hd__dlrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.478500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.680000 0.330000 5.850000 0.665000 ;
        RECT 5.680000 0.665000 6.150000 0.835000 ;
        RECT 5.680000 1.495000 6.065000 1.660000 ;
        RECT 5.680000 1.660000 5.930000 2.465000 ;
        RECT 5.790000 0.835000 6.150000 0.885000 ;
        RECT 5.790000 0.885000 6.360000 1.325000 ;
        RECT 5.790000 1.325000 6.065000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.515000 0.255000 7.765000 0.825000 ;
        RECT 7.515000 1.605000 7.765000 2.465000 ;
        RECT 7.595000 0.825000 7.765000 1.055000 ;
        RECT 7.595000 1.055000 8.195000 1.325000 ;
        RECT 7.595000 1.325000 7.765000 1.605000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.400000 0.995000 5.150000 1.325000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.635000 ;
      RECT 0.085000  0.635000 0.780000 0.805000 ;
      RECT 0.085000  1.795000 0.780000 1.965000 ;
      RECT 0.085000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.455000  1.495000 2.140000 1.665000 ;
      RECT 1.455000  1.665000 1.785000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.140000 0.765000 ;
      RECT 1.535000  0.765000 2.340000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.955000  1.835000 2.270000 2.635000 ;
      RECT 1.970000  0.785000 2.340000 1.095000 ;
      RECT 1.970000  1.095000 2.140000 1.495000 ;
      RECT 2.470000  1.355000 2.755000 1.685000 ;
      RECT 2.715000  0.705000 3.095000 1.035000 ;
      RECT 2.745000  2.255000 3.585000 2.425000 ;
      RECT 2.770000  0.365000 3.500000 0.535000 ;
      RECT 2.925000  1.035000 3.095000 1.575000 ;
      RECT 2.925000  1.575000 3.265000 1.905000 ;
      RECT 2.925000  1.905000 3.125000 1.995000 ;
      RECT 3.270000  2.125000 3.585000 2.255000 ;
      RECT 3.305000  2.075000 3.585000 2.125000 ;
      RECT 3.330000  0.535000 3.500000 0.995000 ;
      RECT 3.330000  0.995000 4.200000 1.165000 ;
      RECT 3.395000  2.015000 3.605000 2.045000 ;
      RECT 3.395000  2.045000 3.585000 2.075000 ;
      RECT 3.415000  1.990000 3.605000 2.015000 ;
      RECT 3.420000  1.975000 3.605000 1.990000 ;
      RECT 3.430000  1.960000 3.605000 1.975000 ;
      RECT 3.435000  1.165000 4.200000 1.325000 ;
      RECT 3.435000  1.325000 3.605000 1.960000 ;
      RECT 3.740000  0.085000 4.070000 0.530000 ;
      RECT 3.755000  2.135000 4.600000 2.635000 ;
      RECT 3.840000  1.535000 5.510000 1.705000 ;
      RECT 3.840000  1.705000 4.940000 1.865000 ;
      RECT 4.270000  0.415000 4.570000 0.655000 ;
      RECT 4.270000  0.655000 5.510000 0.825000 ;
      RECT 4.770000  1.865000 4.940000 2.435000 ;
      RECT 5.110000  0.085000 5.490000 0.485000 ;
      RECT 5.110000  1.875000 5.490000 2.635000 ;
      RECT 5.320000  0.825000 5.510000 0.995000 ;
      RECT 5.320000  0.995000 5.620000 1.325000 ;
      RECT 5.320000  1.325000 5.510000 1.535000 ;
      RECT 6.020000  0.085000 6.360000 0.465000 ;
      RECT 6.100000  1.830000 6.360000 2.635000 ;
      RECT 6.535000  0.255000 6.865000 0.995000 ;
      RECT 6.535000  0.995000 7.425000 1.325000 ;
      RECT 6.535000  1.325000 6.870000 2.465000 ;
      RECT 7.035000  0.085000 7.340000 0.545000 ;
      RECT 7.045000  1.835000 7.340000 2.635000 ;
      RECT 7.935000  0.085000 8.195000 0.885000 ;
      RECT 7.935000  1.495000 8.195000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.445000 2.640000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  1.785000 3.100000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 2.700000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 3.160000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.415000 2.700000 1.460000 ;
      RECT 2.410000 1.600000 2.700000 1.645000 ;
      RECT 2.870000 1.755000 3.160000 1.800000 ;
      RECT 2.870000 1.940000 3.160000 1.985000 ;
  END
END sky130_fd_sc_hd__dlrbp_2
MACRO sky130_fd_sc_hd__dlrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.095000 0.415000 6.355000 2.455000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.500000 0.995000 5.435000 1.325000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.455000  1.495000 2.140000 1.665000 ;
      RECT 1.455000  1.665000 1.785000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.140000 0.765000 ;
      RECT 1.535000  0.765000 2.340000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.955000  1.835000 2.270000 2.635000 ;
      RECT 1.970000  0.785000 2.340000 1.095000 ;
      RECT 1.970000  1.095000 2.140000 1.495000 ;
      RECT 2.470000  1.355000 2.755000 2.005000 ;
      RECT 2.715000  0.705000 3.095000 1.035000 ;
      RECT 2.840000  0.365000 3.500000 0.535000 ;
      RECT 2.900000  2.255000 3.650000 2.425000 ;
      RECT 2.925000  1.035000 3.095000 1.415000 ;
      RECT 2.925000  1.415000 3.265000 1.995000 ;
      RECT 3.330000  0.535000 3.500000 1.025000 ;
      RECT 3.330000  1.025000 4.330000 1.245000 ;
      RECT 3.480000  1.245000 4.330000 1.325000 ;
      RECT 3.480000  1.325000 3.650000 2.255000 ;
      RECT 3.740000  0.085000 4.070000 0.530000 ;
      RECT 3.820000  1.535000 5.925000 1.865000 ;
      RECT 3.820000  2.135000 4.110000 2.635000 ;
      RECT 4.240000  0.255000 4.590000 0.655000 ;
      RECT 4.240000  0.655000 5.925000 0.825000 ;
      RECT 4.300000  2.135000 4.580000 2.635000 ;
      RECT 4.750000  1.865000 4.940000 2.465000 ;
      RECT 5.095000  0.085000 5.925000 0.485000 ;
      RECT 5.110000  2.135000 5.925000 2.635000 ;
      RECT 5.605000  0.825000 5.925000 1.535000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.785000 2.640000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  1.445000 3.100000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.160000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.700000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.755000 2.700000 1.800000 ;
      RECT 2.410000 1.940000 2.700000 1.985000 ;
      RECT 2.870000 1.415000 3.160000 1.460000 ;
      RECT 2.870000 1.600000 3.160000 1.645000 ;
  END
END sky130_fd_sc_hd__dlrtn_1
MACRO sky130_fd_sc_hd__dlrtn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.480500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.595000 0.255000 5.925000 0.485000 ;
        RECT 5.655000 1.875000 5.925000 2.465000 ;
        RECT 5.755000 0.485000 5.925000 0.765000 ;
        RECT 5.755000 0.765000 6.355000 0.865000 ;
        RECT 5.755000 1.425000 6.355000 1.500000 ;
        RECT 5.755000 1.500000 5.925000 1.875000 ;
        RECT 5.760000 1.415000 6.355000 1.425000 ;
        RECT 5.765000 1.410000 6.355000 1.415000 ;
        RECT 5.770000 0.865000 6.355000 0.890000 ;
        RECT 5.775000 1.385000 6.355000 1.410000 ;
        RECT 5.785000 0.890000 6.355000 1.385000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.480000 0.995000 5.170000 1.325000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.455000  1.495000 2.140000 1.665000 ;
      RECT 1.455000  1.665000 1.785000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.140000 0.765000 ;
      RECT 1.535000  0.765000 2.340000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.955000  1.835000 2.270000 2.635000 ;
      RECT 1.960000  0.785000 2.340000 1.095000 ;
      RECT 1.960000  1.095000 2.140000 1.495000 ;
      RECT 2.470000  1.355000 2.755000 2.005000 ;
      RECT 2.675000  0.705000 3.095000 1.145000 ;
      RECT 2.775000  2.255000 3.605000 2.425000 ;
      RECT 2.810000  0.365000 3.500000 0.535000 ;
      RECT 2.925000  1.145000 3.095000 1.415000 ;
      RECT 2.925000  1.415000 3.265000 1.995000 ;
      RECT 3.330000  0.535000 3.500000 1.025000 ;
      RECT 3.330000  1.025000 4.310000 1.245000 ;
      RECT 3.435000  1.245000 4.310000 1.325000 ;
      RECT 3.435000  1.325000 3.605000 2.255000 ;
      RECT 3.735000  0.085000 4.070000 0.530000 ;
      RECT 3.800000  2.135000 4.110000 2.635000 ;
      RECT 3.820000  1.535000 5.585000 1.705000 ;
      RECT 3.820000  1.705000 4.920000 1.865000 ;
      RECT 4.240000  0.255000 4.590000 0.655000 ;
      RECT 4.240000  0.655000 5.585000 0.825000 ;
      RECT 4.280000  2.135000 4.560000 2.635000 ;
      RECT 4.730000  1.865000 4.920000 2.465000 ;
      RECT 5.090000  1.875000 5.460000 2.635000 ;
      RECT 5.095000  0.085000 5.425000 0.485000 ;
      RECT 5.350000  0.995000 5.615000 1.325000 ;
      RECT 5.415000  0.825000 5.585000 0.995000 ;
      RECT 5.415000  1.325000 5.585000 1.535000 ;
      RECT 6.095000  0.085000 6.355000 0.595000 ;
      RECT 6.095000  1.670000 6.355000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.785000 2.640000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  1.445000 3.100000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.160000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.700000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.755000 2.700000 1.800000 ;
      RECT 2.410000 1.940000 2.700000 1.985000 ;
      RECT 2.870000 1.415000 3.160000 1.460000 ;
      RECT 2.870000 1.600000 3.160000 1.645000 ;
  END
END sky130_fd_sc_hd__dlrtn_2
MACRO sky130_fd_sc_hd__dlrtn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 0.955000 1.795000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.014750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.610000 0.255000 5.965000 0.485000 ;
        RECT 5.680000 1.875000 5.965000 2.465000 ;
        RECT 5.795000 0.485000 5.965000 0.765000 ;
        RECT 5.795000 0.765000 7.275000 1.325000 ;
        RECT 5.795000 1.325000 5.965000 1.875000 ;
        RECT 6.575000 0.255000 6.775000 0.765000 ;
        RECT 6.575000 1.325000 6.775000 2.465000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.505000 0.995000 5.145000 1.325000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.360000 2.805000 ;
        RECT 0.515000 2.135000 0.845000 2.635000 ;
        RECT 1.960000 1.835000 2.275000 2.635000 ;
        RECT 3.825000 2.135000 4.115000 2.635000 ;
        RECT 4.305000 2.135000 4.585000 2.635000 ;
        RECT 5.115000 1.875000 5.485000 2.635000 ;
        RECT 6.135000 1.495000 6.405000 2.635000 ;
        RECT 6.945000 1.495000 7.275000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.460000  1.495000 2.145000 1.665000 ;
      RECT 1.460000  1.665000 1.790000 2.415000 ;
      RECT 1.540000  0.345000 1.710000 0.615000 ;
      RECT 1.540000  0.615000 2.145000 0.765000 ;
      RECT 1.540000  0.765000 2.345000 0.785000 ;
      RECT 1.880000  0.085000 2.210000 0.445000 ;
      RECT 1.975000  0.785000 2.345000 1.095000 ;
      RECT 1.975000  1.095000 2.145000 1.495000 ;
      RECT 2.475000  1.355000 2.760000 2.005000 ;
      RECT 2.720000  0.705000 3.100000 1.035000 ;
      RECT 2.845000  0.365000 3.505000 0.535000 ;
      RECT 2.905000  2.255000 3.655000 2.425000 ;
      RECT 2.930000  1.035000 3.100000 1.415000 ;
      RECT 2.930000  1.415000 3.270000 1.995000 ;
      RECT 3.335000  0.535000 3.505000 1.025000 ;
      RECT 3.335000  1.025000 4.315000 1.245000 ;
      RECT 3.485000  1.245000 4.315000 1.325000 ;
      RECT 3.485000  1.325000 3.655000 2.255000 ;
      RECT 3.745000  0.085000 4.075000 0.530000 ;
      RECT 3.825000  1.535000 5.625000 1.705000 ;
      RECT 3.825000  1.705000 4.945000 1.865000 ;
      RECT 4.245000  0.255000 4.595000 0.655000 ;
      RECT 4.245000  0.655000 5.625000 0.825000 ;
      RECT 4.755000  1.865000 4.945000 2.465000 ;
      RECT 5.100000  0.085000 5.440000 0.485000 ;
      RECT 5.455000  0.825000 5.625000 1.535000 ;
      RECT 6.135000  0.085000 6.405000 0.595000 ;
      RECT 6.945000  0.085000 7.275000 0.595000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.475000  1.785000 2.645000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.935000  1.445000 3.105000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.165000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.705000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.415000 1.755000 2.705000 1.800000 ;
      RECT 2.415000 1.940000 2.705000 1.985000 ;
      RECT 2.875000 1.415000 3.165000 1.460000 ;
      RECT 2.875000 1.600000 3.165000 1.645000 ;
  END
END sky130_fd_sc_hd__dlrtn_4
MACRO sky130_fd_sc_hd__dlrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.955000 1.765000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.610000 0.345000 5.895000 0.745000 ;
        RECT 5.635000 1.670000 5.895000 2.455000 ;
        RECT 5.725000 0.745000 5.895000 1.670000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.745000 0.345000 4.975000 0.995000 ;
        RECT 4.745000 0.995000 5.075000 1.325000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.325000 1.625000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  1.795000 0.775000 1.965000 ;
      RECT 0.085000  1.965000 0.345000 2.465000 ;
      RECT 0.170000  0.345000 0.345000 0.635000 ;
      RECT 0.170000  0.635000 0.775000 0.805000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.605000  0.805000 0.775000 1.070000 ;
      RECT 0.605000  1.070000 0.835000 1.400000 ;
      RECT 0.605000  1.400000 0.775000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.235000 2.465000 ;
      RECT 1.430000  1.495000 2.115000 1.665000 ;
      RECT 1.430000  1.665000 1.785000 2.415000 ;
      RECT 1.510000  0.345000 1.705000 0.615000 ;
      RECT 1.510000  0.615000 2.115000 0.765000 ;
      RECT 1.510000  0.765000 2.335000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.945000  0.785000 2.335000 1.095000 ;
      RECT 1.945000  1.095000 2.115000 1.495000 ;
      RECT 1.955000  1.835000 2.245000 2.635000 ;
      RECT 2.445000  1.355000 2.835000 1.625000 ;
      RECT 2.445000  1.625000 2.760000 1.685000 ;
      RECT 2.690000  0.765000 3.245000 1.095000 ;
      RECT 2.810000  2.255000 3.625000 2.425000 ;
      RECT 2.815000  0.365000 3.585000 0.535000 ;
      RECT 2.900000  1.785000 3.265000 1.995000 ;
      RECT 3.005000  1.095000 3.245000 1.635000 ;
      RECT 3.005000  1.635000 3.265000 1.785000 ;
      RECT 3.415000  0.535000 3.585000 0.995000 ;
      RECT 3.415000  0.995000 4.175000 1.165000 ;
      RECT 3.455000  1.165000 4.175000 1.325000 ;
      RECT 3.455000  1.325000 3.625000 2.255000 ;
      RECT 3.755000  0.085000 4.025000 0.610000 ;
      RECT 3.815000  1.535000 5.465000 1.735000 ;
      RECT 3.815000  1.735000 4.965000 1.865000 ;
      RECT 3.930000  2.135000 4.445000 2.635000 ;
      RECT 4.195000  0.295000 4.575000 0.805000 ;
      RECT 4.345000  0.805000 4.575000 1.505000 ;
      RECT 4.345000  1.505000 5.465000 1.535000 ;
      RECT 4.625000  1.865000 4.965000 2.435000 ;
      RECT 5.135000  1.915000 5.465000 2.635000 ;
      RECT 5.155000  0.085000 5.440000 0.715000 ;
      RECT 5.245000  0.995000 5.555000 1.325000 ;
      RECT 5.245000  1.325000 5.465000 1.505000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  1.445000 0.775000 1.615000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  1.785000 1.235000 1.955000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  1.445000 2.615000 1.615000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.925000  1.785000 3.095000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 0.545000 1.415000 0.835000 1.460000 ;
      RECT 0.545000 1.460000 2.675000 1.600000 ;
      RECT 0.545000 1.600000 0.835000 1.645000 ;
      RECT 1.005000 1.755000 1.295000 1.800000 ;
      RECT 1.005000 1.800000 3.155000 1.940000 ;
      RECT 1.005000 1.940000 1.295000 1.985000 ;
      RECT 2.385000 1.415000 2.675000 1.460000 ;
      RECT 2.385000 1.600000 2.675000 1.645000 ;
      RECT 2.865000 1.755000 3.155000 1.800000 ;
      RECT 2.865000 1.940000 3.155000 1.985000 ;
  END
END sky130_fd_sc_hd__dlrtp_1
MACRO sky130_fd_sc_hd__dlrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.440000 0.955000 1.770000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.480500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.595000 0.255000 5.925000 0.485000 ;
        RECT 5.655000 1.875000 5.925000 2.465000 ;
        RECT 5.755000 0.485000 5.925000 0.765000 ;
        RECT 5.755000 0.765000 6.355000 0.865000 ;
        RECT 5.755000 1.425000 6.355000 1.500000 ;
        RECT 5.755000 1.500000 5.925000 1.875000 ;
        RECT 5.760000 1.415000 6.355000 1.425000 ;
        RECT 5.765000 1.410000 6.355000 1.415000 ;
        RECT 5.770000 0.865000 6.355000 0.890000 ;
        RECT 5.775000 1.385000 6.355000 1.410000 ;
        RECT 5.785000 0.890000 6.355000 1.385000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.480000 0.995000 4.815000 1.035000 ;
        RECT 4.480000 1.035000 5.240000 1.325000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.985000 0.330000 1.625000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.635000 ;
      RECT 0.085000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.435000  1.495000 2.120000 1.665000 ;
      RECT 1.435000  1.665000 1.785000 2.415000 ;
      RECT 1.515000  0.345000 1.705000 0.615000 ;
      RECT 1.515000  0.615000 2.120000 0.765000 ;
      RECT 1.515000  0.765000 2.335000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.950000  0.785000 2.335000 1.095000 ;
      RECT 1.950000  1.095000 2.120000 1.495000 ;
      RECT 1.955000  1.835000 2.250000 2.635000 ;
      RECT 2.450000  1.355000 2.755000 1.685000 ;
      RECT 2.585000  0.735000 3.100000 1.040000 ;
      RECT 2.770000  0.365000 3.445000 0.535000 ;
      RECT 2.770000  2.255000 3.580000 2.425000 ;
      RECT 2.905000  1.780000 3.265000 1.910000 ;
      RECT 2.905000  1.910000 3.175000 1.995000 ;
      RECT 2.930000  1.040000 3.100000 1.570000 ;
      RECT 2.930000  1.570000 3.265000 1.780000 ;
      RECT 3.270000  0.535000 3.445000 0.995000 ;
      RECT 3.270000  0.995000 4.220000 1.325000 ;
      RECT 3.410000  2.000000 3.605000 2.085000 ;
      RECT 3.410000  2.085000 3.580000 2.255000 ;
      RECT 3.415000  1.995000 3.605000 2.000000 ;
      RECT 3.420000  1.985000 3.605000 1.995000 ;
      RECT 3.435000  1.325000 3.605000 1.985000 ;
      RECT 3.720000  0.085000 4.060000 0.530000 ;
      RECT 3.750000  2.175000 4.090000 2.635000 ;
      RECT 3.775000  1.535000 5.585000 1.705000 ;
      RECT 3.775000  1.705000 4.970000 1.865000 ;
      RECT 4.240000  0.255000 4.580000 0.655000 ;
      RECT 4.240000  0.655000 5.095000 0.695000 ;
      RECT 4.240000  0.695000 5.585000 0.825000 ;
      RECT 4.280000  2.135000 4.560000 2.635000 ;
      RECT 4.800000  1.865000 4.970000 2.465000 ;
      RECT 4.955000  0.825000 5.585000 0.865000 ;
      RECT 5.140000  1.875000 5.485000 2.635000 ;
      RECT 5.255000  0.085000 5.425000 0.525000 ;
      RECT 5.415000  0.865000 5.585000 0.995000 ;
      RECT 5.415000  0.995000 5.615000 1.325000 ;
      RECT 5.415000  1.325000 5.585000 1.535000 ;
      RECT 6.095000  0.085000 6.355000 0.595000 ;
      RECT 6.095000  1.670000 6.355000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.450000  1.445000 2.620000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.925000  1.785000 3.095000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 2.680000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 3.155000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.390000 1.415000 2.680000 1.460000 ;
      RECT 2.390000 1.600000 2.680000 1.645000 ;
      RECT 2.865000 1.755000 3.155000 1.800000 ;
      RECT 2.865000 1.940000 3.155000 1.985000 ;
  END
END sky130_fd_sc_hd__dlrtp_2
MACRO sky130_fd_sc_hd__dlrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 0.955000 1.795000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.014750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.610000 0.255000 5.965000 0.485000 ;
        RECT 5.680000 1.875000 5.965000 2.465000 ;
        RECT 5.795000 0.485000 5.965000 0.765000 ;
        RECT 5.795000 0.765000 7.275000 1.325000 ;
        RECT 5.795000 1.325000 5.965000 1.875000 ;
        RECT 6.575000 0.255000 6.775000 0.765000 ;
        RECT 6.575000 1.325000 6.775000 2.465000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.505000 0.995000 5.145000 1.325000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.360000 2.805000 ;
        RECT 0.515000 2.135000 0.845000 2.635000 ;
        RECT 1.960000 1.835000 2.275000 2.635000 ;
        RECT 3.825000 2.135000 4.115000 2.635000 ;
        RECT 4.305000 2.135000 4.585000 2.635000 ;
        RECT 5.115000 1.875000 5.485000 2.635000 ;
        RECT 6.135000 1.495000 6.405000 2.635000 ;
        RECT 6.945000 1.495000 7.275000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.460000  1.495000 2.145000 1.665000 ;
      RECT 1.460000  1.665000 1.790000 2.415000 ;
      RECT 1.540000  0.345000 1.710000 0.615000 ;
      RECT 1.540000  0.615000 2.145000 0.765000 ;
      RECT 1.540000  0.765000 2.345000 0.785000 ;
      RECT 1.880000  0.085000 2.210000 0.445000 ;
      RECT 1.975000  0.785000 2.345000 1.095000 ;
      RECT 1.975000  1.095000 2.145000 1.495000 ;
      RECT 2.475000  1.355000 2.760000 1.685000 ;
      RECT 2.720000  0.705000 3.100000 1.035000 ;
      RECT 2.845000  0.365000 3.505000 0.535000 ;
      RECT 2.905000  2.255000 3.655000 2.425000 ;
      RECT 2.930000  1.035000 3.100000 1.575000 ;
      RECT 2.930000  1.575000 3.270000 1.995000 ;
      RECT 3.335000  0.535000 3.505000 0.995000 ;
      RECT 3.335000  0.995000 4.235000 1.165000 ;
      RECT 3.485000  1.165000 4.235000 1.325000 ;
      RECT 3.485000  1.325000 3.655000 2.255000 ;
      RECT 3.745000  0.085000 4.075000 0.530000 ;
      RECT 3.825000  1.535000 5.625000 1.705000 ;
      RECT 3.825000  1.705000 4.945000 1.865000 ;
      RECT 4.265000  0.255000 4.595000 0.655000 ;
      RECT 4.265000  0.655000 5.625000 0.825000 ;
      RECT 4.755000  1.865000 4.945000 2.465000 ;
      RECT 5.100000  0.085000 5.440000 0.485000 ;
      RECT 5.455000  0.825000 5.625000 1.535000 ;
      RECT 6.135000  0.085000 6.405000 0.595000 ;
      RECT 6.945000  0.085000 7.275000 0.595000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.475000  1.445000 2.645000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.935000  1.785000 3.105000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 2.705000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 3.165000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.415000 1.415000 2.705000 1.460000 ;
      RECT 2.415000 1.600000 2.705000 1.645000 ;
      RECT 2.875000 1.755000 3.165000 1.800000 ;
      RECT 2.875000 1.940000 3.165000 1.985000 ;
  END
END sky130_fd_sc_hd__dlrtp_4
MACRO sky130_fd_sc_hd__dlxbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445000 0.955000 1.785000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.140000 0.415000 5.480000 0.745000 ;
        RECT 5.140000 1.670000 5.480000 2.465000 ;
        RECT 5.310000 0.745000 5.480000 1.670000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.555000 0.255000 6.815000 0.825000 ;
        RECT 6.555000 1.505000 6.815000 2.465000 ;
        RECT 6.625000 0.825000 6.815000 1.505000 ;
    END
  END Q_N
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.090000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.480000  1.495000 2.165000 1.665000 ;
      RECT 1.480000  1.665000 1.810000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.165000 0.785000 ;
      RECT 1.875000  0.085000 2.230000 0.445000 ;
      RECT 1.980000  1.835000 2.295000 2.635000 ;
      RECT 1.995000  0.785000 2.165000 0.905000 ;
      RECT 1.995000  0.905000 2.365000 1.235000 ;
      RECT 1.995000  1.235000 2.165000 1.495000 ;
      RECT 2.495000  1.355000 2.780000 2.005000 ;
      RECT 2.565000  0.705000 3.120000 1.035000 ;
      RECT 2.790000  0.365000 3.525000 0.535000 ;
      RECT 2.920000  2.105000 3.620000 2.115000 ;
      RECT 2.920000  2.115000 3.615000 2.130000 ;
      RECT 2.920000  2.130000 3.610000 2.275000 ;
      RECT 2.950000  1.035000 3.120000 1.415000 ;
      RECT 2.950000  1.415000 3.290000 1.910000 ;
      RECT 3.355000  0.535000 3.525000 0.995000 ;
      RECT 3.355000  0.995000 4.225000 1.165000 ;
      RECT 3.360000  2.075000 3.630000 2.090000 ;
      RECT 3.360000  2.090000 3.625000 2.105000 ;
      RECT 3.375000  2.060000 3.630000 2.075000 ;
      RECT 3.420000  2.030000 3.630000 2.060000 ;
      RECT 3.430000  2.015000 3.630000 2.030000 ;
      RECT 3.460000  1.165000 4.225000 1.325000 ;
      RECT 3.460000  1.325000 3.630000 2.015000 ;
      RECT 3.765000  0.085000 4.095000 0.610000 ;
      RECT 3.780000  2.175000 3.950000 2.635000 ;
      RECT 3.800000  1.535000 4.580000 1.620000 ;
      RECT 3.800000  1.620000 4.550000 1.865000 ;
      RECT 4.300000  0.415000 4.470000 0.660000 ;
      RECT 4.300000  0.660000 4.580000 0.840000 ;
      RECT 4.300000  1.865000 4.550000 2.435000 ;
      RECT 4.395000  0.840000 4.580000 0.995000 ;
      RECT 4.395000  0.995000 5.140000 1.325000 ;
      RECT 4.395000  1.325000 4.580000 1.535000 ;
      RECT 4.640000  0.085000 4.970000 0.495000 ;
      RECT 4.720000  1.830000 4.970000 2.635000 ;
      RECT 5.660000  0.255000 5.910000 0.995000 ;
      RECT 5.660000  0.995000 6.455000 1.325000 ;
      RECT 5.660000  1.325000 5.910000 2.465000 ;
      RECT 6.090000  0.085000 6.385000 0.545000 ;
      RECT 6.090000  1.835000 6.385000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.495000  1.785000 2.665000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.955000  1.445000 3.125000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.185000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.725000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.435000 1.755000 2.725000 1.800000 ;
      RECT 2.435000 1.940000 2.725000 1.985000 ;
      RECT 2.895000 1.415000 3.185000 1.460000 ;
      RECT 2.895000 1.600000 3.185000 1.645000 ;
  END
END sky130_fd_sc_hd__dlxbn_1
MACRO sky130_fd_sc_hd__dlxbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxbn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 0.955000 1.810000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.215000 0.415000 5.465000 0.660000 ;
        RECT 5.215000 0.660000 5.500000 0.825000 ;
        RECT 5.215000 1.495000 5.500000 1.710000 ;
        RECT 5.215000 1.710000 5.465000 2.455000 ;
        RECT 5.330000 0.825000 5.500000 0.995000 ;
        RECT 5.330000 0.995000 5.905000 1.325000 ;
        RECT 5.330000 1.325000 5.500000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.050000 0.255000 7.305000 0.825000 ;
        RECT 7.050000 1.445000 7.305000 2.465000 ;
        RECT 7.095000 0.825000 7.305000 1.055000 ;
        RECT 7.095000 1.055000 7.735000 1.325000 ;
        RECT 7.095000 1.325000 7.305000 1.445000 ;
    END
  END Q_N
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.475000  1.495000 2.160000 1.665000 ;
      RECT 1.475000  1.665000 1.805000 2.415000 ;
      RECT 1.555000  0.345000 1.725000 0.615000 ;
      RECT 1.555000  0.615000 2.160000 0.765000 ;
      RECT 1.555000  0.765000 2.360000 0.785000 ;
      RECT 1.895000  0.085000 2.225000 0.445000 ;
      RECT 1.975000  1.835000 2.290000 2.635000 ;
      RECT 1.990000  0.785000 2.360000 1.095000 ;
      RECT 1.990000  1.095000 2.160000 1.495000 ;
      RECT 2.490000  1.355000 2.775000 2.005000 ;
      RECT 2.735000  0.705000 3.115000 1.035000 ;
      RECT 2.860000  0.365000 3.520000 0.535000 ;
      RECT 2.920000  2.255000 3.670000 2.425000 ;
      RECT 2.945000  1.035000 3.115000 1.415000 ;
      RECT 2.945000  1.415000 3.285000 1.995000 ;
      RECT 3.350000  0.535000 3.520000 0.995000 ;
      RECT 3.350000  0.995000 4.220000 1.165000 ;
      RECT 3.500000  1.165000 4.220000 1.325000 ;
      RECT 3.500000  1.325000 3.670000 2.255000 ;
      RECT 3.760000  0.085000 4.090000 0.825000 ;
      RECT 3.840000  2.135000 4.140000 2.635000 ;
      RECT 3.860000  1.535000 4.580000 1.865000 ;
      RECT 4.360000  0.415000 4.580000 0.825000 ;
      RECT 4.360000  1.865000 4.580000 2.435000 ;
      RECT 4.410000  0.825000 4.580000 0.995000 ;
      RECT 4.410000  0.995000 5.160000 1.325000 ;
      RECT 4.410000  1.325000 4.580000 1.535000 ;
      RECT 4.760000  0.085000 5.045000 0.825000 ;
      RECT 4.760000  1.495000 5.045000 2.635000 ;
      RECT 5.635000  0.085000 5.905000 0.545000 ;
      RECT 5.635000  1.835000 5.905000 2.635000 ;
      RECT 6.075000  0.255000 6.405000 0.995000 ;
      RECT 6.075000  0.995000 6.925000 1.325000 ;
      RECT 6.075000  1.325000 6.405000 2.465000 ;
      RECT 6.585000  0.085000 6.880000 0.545000 ;
      RECT 6.585000  1.835000 6.880000 2.635000 ;
      RECT 7.475000  0.085000 7.735000 0.885000 ;
      RECT 7.475000  1.495000 7.735000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.490000  1.785000 2.660000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.950000  1.445000 3.120000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.180000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.720000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.430000 1.755000 2.720000 1.800000 ;
      RECT 2.430000 1.940000 2.720000 1.985000 ;
      RECT 2.890000 1.415000 3.180000 1.460000 ;
      RECT 2.890000 1.600000 3.180000 1.645000 ;
  END
END sky130_fd_sc_hd__dlxbn_2
MACRO sky130_fd_sc_hd__dlxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 0.955000 1.685000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.140000 0.255000 5.490000 0.820000 ;
        RECT 5.140000 1.670000 5.490000 2.455000 ;
        RECT 5.320000 0.820000 5.490000 1.670000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.555000 0.255000 6.815000 0.825000 ;
        RECT 6.555000 1.445000 6.815000 2.465000 ;
        RECT 6.600000 0.825000 6.815000 1.445000 ;
    END
  END Q_N
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.090000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.430000  1.495000 2.115000 1.665000 ;
      RECT 1.430000  1.665000 1.795000 2.415000 ;
      RECT 1.510000  0.345000 1.705000 0.615000 ;
      RECT 1.510000  0.615000 2.135000 0.785000 ;
      RECT 1.855000  0.785000 2.135000 0.875000 ;
      RECT 1.855000  0.875000 2.335000 1.235000 ;
      RECT 1.855000  1.235000 2.115000 1.495000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.965000  1.835000 2.245000 2.635000 ;
      RECT 2.465000  1.355000 2.795000 1.685000 ;
      RECT 2.580000  0.705000 3.135000 1.065000 ;
      RECT 2.750000  2.255000 3.610000 2.425000 ;
      RECT 2.800000  0.365000 3.475000 0.535000 ;
      RECT 2.965000  1.065000 3.135000 1.575000 ;
      RECT 2.965000  1.575000 3.290000 1.910000 ;
      RECT 2.965000  1.910000 3.195000 1.995000 ;
      RECT 3.305000  0.535000 3.475000 0.995000 ;
      RECT 3.305000  0.995000 4.175000 1.165000 ;
      RECT 3.425000  2.035000 3.650000 2.065000 ;
      RECT 3.425000  2.065000 3.630000 2.090000 ;
      RECT 3.425000  2.090000 3.610000 2.255000 ;
      RECT 3.430000  2.020000 3.650000 2.035000 ;
      RECT 3.435000  2.010000 3.650000 2.020000 ;
      RECT 3.440000  1.995000 3.650000 2.010000 ;
      RECT 3.460000  1.165000 4.175000 1.325000 ;
      RECT 3.460000  1.325000 3.650000 1.995000 ;
      RECT 3.700000  0.085000 4.045000 0.530000 ;
      RECT 3.780000  2.175000 3.980000 2.635000 ;
      RECT 3.820000  1.535000 4.515000 1.865000 ;
      RECT 4.285000  0.415000 4.550000 0.745000 ;
      RECT 4.285000  1.865000 4.515000 2.435000 ;
      RECT 4.345000  0.745000 4.550000 0.995000 ;
      RECT 4.345000  0.995000 5.150000 1.325000 ;
      RECT 4.345000  1.325000 4.515000 1.535000 ;
      RECT 4.685000  1.570000 4.970000 2.635000 ;
      RECT 4.720000  0.085000 4.970000 0.715000 ;
      RECT 5.660000  0.255000 5.910000 0.995000 ;
      RECT 5.660000  0.995000 6.430000 1.325000 ;
      RECT 5.660000  1.325000 5.910000 2.465000 ;
      RECT 6.090000  0.085000 6.385000 0.545000 ;
      RECT 6.090000  1.835000 6.385000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.555000  1.445000 2.725000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.965000  1.785000 3.135000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 2.785000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 3.195000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.495000 1.415000 2.785000 1.460000 ;
      RECT 2.495000 1.600000 2.785000 1.645000 ;
      RECT 2.905000 1.755000 3.195000 1.800000 ;
      RECT 2.905000 1.940000 3.195000 1.985000 ;
  END
END sky130_fd_sc_hd__dlxbp_1
MACRO sky130_fd_sc_hd__dlxtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.955000 1.765000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.175000 0.415000 5.435000 0.745000 ;
        RECT 5.175000 1.670000 5.435000 2.455000 ;
        RECT 5.265000 0.745000 5.435000 1.670000 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.430000  1.495000 2.115000 1.665000 ;
      RECT 1.430000  1.665000 1.785000 2.415000 ;
      RECT 1.510000  0.345000 1.705000 0.615000 ;
      RECT 1.510000  0.615000 2.115000 0.765000 ;
      RECT 1.510000  0.765000 2.320000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.945000  0.785000 2.320000 1.235000 ;
      RECT 1.945000  1.235000 2.115000 1.495000 ;
      RECT 1.955000  1.835000 2.245000 2.635000 ;
      RECT 2.445000  1.355000 2.780000 2.005000 ;
      RECT 2.560000  0.735000 3.265000 1.040000 ;
      RECT 2.745000  2.255000 3.605000 2.425000 ;
      RECT 2.765000  0.365000 3.605000 0.535000 ;
      RECT 2.950000  1.040000 3.265000 1.560000 ;
      RECT 2.950000  1.560000 3.285000 1.910000 ;
      RECT 3.295000  2.090000 3.620000 2.105000 ;
      RECT 3.295000  2.105000 3.605000 2.255000 ;
      RECT 3.390000  2.045000 3.645000 2.065000 ;
      RECT 3.390000  2.065000 3.630000 2.085000 ;
      RECT 3.390000  2.085000 3.620000 2.090000 ;
      RECT 3.405000  2.035000 3.645000 2.045000 ;
      RECT 3.430000  2.010000 3.645000 2.035000 ;
      RECT 3.435000  0.535000 3.605000 0.995000 ;
      RECT 3.435000  0.995000 4.200000 1.325000 ;
      RECT 3.435000  1.325000 3.645000 1.450000 ;
      RECT 3.455000  1.450000 3.645000 2.010000 ;
      RECT 3.775000  0.085000 4.045000 0.545000 ;
      RECT 3.775000  2.175000 4.095000 2.635000 ;
      RECT 3.815000  1.535000 4.540000 1.865000 ;
      RECT 4.295000  0.260000 4.540000 0.720000 ;
      RECT 4.295000  1.865000 4.540000 2.435000 ;
      RECT 4.370000  0.720000 4.540000 0.995000 ;
      RECT 4.370000  0.995000 5.095000 1.325000 ;
      RECT 4.370000  1.325000 4.540000 1.535000 ;
      RECT 4.720000  1.570000 5.005000 2.635000 ;
      RECT 4.755000  0.085000 4.980000 0.715000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  1.785000 2.615000 1.955000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.950000  1.445000 3.120000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.180000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.675000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.385000 1.755000 2.675000 1.800000 ;
      RECT 2.385000 1.940000 2.675000 1.985000 ;
      RECT 2.890000 1.415000 3.180000 1.460000 ;
      RECT 2.890000 1.600000 3.180000 1.645000 ;
  END
END sky130_fd_sc_hd__dlxtn_1
MACRO sky130_fd_sc_hd__dlxtn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxtn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 0.955000 1.810000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.215000 0.415000 5.465000 0.685000 ;
        RECT 5.215000 0.685000 5.500000 0.825000 ;
        RECT 5.215000 1.495000 5.500000 1.640000 ;
        RECT 5.215000 1.640000 5.465000 2.455000 ;
        RECT 5.330000 0.825000 5.500000 0.995000 ;
        RECT 5.330000 0.995000 5.895000 1.325000 ;
        RECT 5.330000 1.325000 5.500000 1.495000 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.475000  1.495000 2.160000 1.665000 ;
      RECT 1.475000  1.665000 1.805000 2.415000 ;
      RECT 1.555000  0.345000 1.725000 0.615000 ;
      RECT 1.555000  0.615000 2.160000 0.765000 ;
      RECT 1.555000  0.765000 2.360000 0.785000 ;
      RECT 1.895000  0.085000 2.225000 0.445000 ;
      RECT 1.975000  1.835000 2.290000 2.635000 ;
      RECT 1.990000  0.785000 2.360000 1.095000 ;
      RECT 1.990000  1.095000 2.160000 1.495000 ;
      RECT 2.490000  1.355000 2.775000 2.005000 ;
      RECT 2.735000  0.705000 3.115000 1.035000 ;
      RECT 2.860000  0.365000 3.520000 0.535000 ;
      RECT 2.920000  2.255000 3.670000 2.425000 ;
      RECT 2.945000  1.035000 3.115000 1.415000 ;
      RECT 2.945000  1.415000 3.285000 1.995000 ;
      RECT 3.350000  0.535000 3.520000 0.995000 ;
      RECT 3.350000  0.995000 4.220000 1.165000 ;
      RECT 3.500000  1.165000 4.220000 1.325000 ;
      RECT 3.500000  1.325000 3.670000 2.255000 ;
      RECT 3.760000  0.085000 4.090000 0.825000 ;
      RECT 3.840000  2.135000 4.140000 2.635000 ;
      RECT 3.860000  1.535000 4.580000 1.865000 ;
      RECT 4.360000  0.415000 4.580000 0.825000 ;
      RECT 4.360000  1.865000 4.580000 2.435000 ;
      RECT 4.410000  0.825000 4.580000 0.995000 ;
      RECT 4.410000  0.995000 5.160000 1.325000 ;
      RECT 4.410000  1.325000 4.580000 1.535000 ;
      RECT 4.760000  0.085000 5.045000 0.825000 ;
      RECT 4.760000  1.495000 5.045000 2.635000 ;
      RECT 5.635000  0.085000 5.895000 0.550000 ;
      RECT 5.635000  1.755000 5.895000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.490000  1.785000 2.660000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.950000  1.445000 3.120000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.180000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.720000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.430000 1.755000 2.720000 1.800000 ;
      RECT 2.430000 1.940000 2.720000 1.985000 ;
      RECT 2.890000 1.415000 3.180000 1.460000 ;
      RECT 2.890000 1.600000 3.180000 1.645000 ;
  END
END sky130_fd_sc_hd__dlxtn_2
MACRO sky130_fd_sc_hd__dlxtn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxtn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.240000 0.415000 5.525000 0.745000 ;
        RECT 5.240000 1.495000 5.525000 2.455000 ;
        RECT 5.355000 0.745000 5.525000 0.995000 ;
        RECT 5.355000 0.995000 6.815000 1.325000 ;
        RECT 5.355000 1.325000 5.525000 1.495000 ;
        RECT 6.115000 0.385000 6.385000 0.995000 ;
        RECT 6.115000 1.325000 6.385000 2.455000 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.090000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.455000  1.495000 2.140000 1.665000 ;
      RECT 1.455000  1.665000 1.785000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.140000 0.765000 ;
      RECT 1.535000  0.765000 2.340000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.955000  1.835000 2.270000 2.635000 ;
      RECT 1.970000  0.785000 2.340000 1.095000 ;
      RECT 1.970000  1.095000 2.140000 1.495000 ;
      RECT 2.470000  1.355000 2.755000 2.005000 ;
      RECT 2.715000  0.705000 3.095000 1.035000 ;
      RECT 2.840000  0.365000 3.500000 0.535000 ;
      RECT 2.900000  2.255000 3.650000 2.425000 ;
      RECT 2.925000  1.035000 3.095000 1.415000 ;
      RECT 2.925000  1.415000 3.265000 1.995000 ;
      RECT 3.330000  0.535000 3.500000 0.995000 ;
      RECT 3.330000  0.995000 4.200000 1.165000 ;
      RECT 3.480000  1.165000 4.200000 1.325000 ;
      RECT 3.480000  1.325000 3.650000 2.255000 ;
      RECT 3.740000  0.085000 4.070000 0.530000 ;
      RECT 3.820000  2.135000 4.120000 2.635000 ;
      RECT 3.840000  1.535000 4.605000 1.865000 ;
      RECT 4.385000  0.415000 4.605000 0.745000 ;
      RECT 4.385000  1.865000 4.605000 2.435000 ;
      RECT 4.435000  0.745000 4.605000 0.995000 ;
      RECT 4.435000  0.995000 5.185000 1.325000 ;
      RECT 4.435000  1.325000 4.605000 1.535000 ;
      RECT 4.785000  0.085000 5.070000 0.715000 ;
      RECT 4.785000  1.495000 5.070000 2.635000 ;
      RECT 5.695000  0.085000 5.945000 0.825000 ;
      RECT 5.695000  1.495000 5.945000 2.635000 ;
      RECT 6.555000  0.085000 6.815000 0.715000 ;
      RECT 6.555000  1.495000 6.815000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.785000 2.640000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  1.445000 3.100000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.160000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.700000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.755000 2.700000 1.800000 ;
      RECT 2.410000 1.940000 2.700000 1.985000 ;
      RECT 2.870000 1.415000 3.160000 1.460000 ;
      RECT 2.870000 1.600000 3.160000 1.645000 ;
  END
END sky130_fd_sc_hd__dlxtn_4
MACRO sky130_fd_sc_hd__dlxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.470250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.150000 0.415000 5.435000 0.745000 ;
        RECT 5.150000 1.670000 5.435000 2.455000 ;
        RECT 5.265000 0.745000 5.435000 1.670000 ;
    END
  END Q
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.985000 0.330000 1.625000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.455000  1.495000 2.140000 1.665000 ;
      RECT 1.455000  1.665000 1.785000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.140000 0.765000 ;
      RECT 1.535000  0.765000 2.340000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.955000  1.835000 2.270000 2.635000 ;
      RECT 1.970000  0.785000 2.340000 1.095000 ;
      RECT 1.970000  1.095000 2.140000 1.495000 ;
      RECT 2.470000  1.355000 2.755000 1.685000 ;
      RECT 2.715000  0.705000 3.095000 1.035000 ;
      RECT 2.770000  2.255000 3.605000 2.425000 ;
      RECT 2.840000  0.365000 3.500000 0.535000 ;
      RECT 2.925000  1.035000 3.095000 1.575000 ;
      RECT 2.925000  1.575000 3.265000 1.995000 ;
      RECT 3.330000  0.535000 3.500000 0.995000 ;
      RECT 3.330000  0.995000 4.175000 1.165000 ;
      RECT 3.435000  1.165000 4.175000 1.325000 ;
      RECT 3.435000  1.325000 3.605000 2.255000 ;
      RECT 3.685000  0.085000 4.015000 0.530000 ;
      RECT 3.775000  2.135000 3.945000 2.635000 ;
      RECT 3.840000  1.535000 4.515000 1.865000 ;
      RECT 4.295000  0.415000 4.515000 0.745000 ;
      RECT 4.295000  1.865000 4.515000 2.435000 ;
      RECT 4.345000  0.745000 4.515000 0.995000 ;
      RECT 4.345000  0.995000 5.095000 1.325000 ;
      RECT 4.345000  1.325000 4.515000 1.535000 ;
      RECT 4.695000  0.085000 4.900000 0.715000 ;
      RECT 4.695000  1.570000 4.900000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.445000 2.640000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  1.785000 3.100000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 2.700000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 3.160000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.415000 2.700000 1.460000 ;
      RECT 2.410000 1.600000 2.700000 1.645000 ;
      RECT 2.870000 1.755000 3.160000 1.800000 ;
      RECT 2.870000 1.940000 3.160000 1.985000 ;
  END
END sky130_fd_sc_hd__dlxtp_1
MACRO sky130_fd_sc_hd__dlygate4sd1_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlygate4sd1_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.555000 1.615000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.410000 0.255000 2.700000 0.825000 ;
        RECT 2.440000 1.495000 2.700000 2.465000 ;
        RECT 2.530000 0.825000 2.700000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.085000 0.310000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  1.785000 0.895000 2.005000 ;
      RECT 0.085000  2.005000 0.380000 2.465000 ;
      RECT 0.095000  0.255000 0.380000 0.715000 ;
      RECT 0.095000  0.715000 0.895000 0.885000 ;
      RECT 0.550000  0.085000 0.765000 0.545000 ;
      RECT 0.550000  2.175000 0.765000 2.635000 ;
      RECT 0.725000  0.885000 0.895000 0.995000 ;
      RECT 0.725000  0.995000 0.980000 1.325000 ;
      RECT 0.725000  1.325000 0.895000 1.785000 ;
      RECT 0.935000  0.255000 1.320000 0.545000 ;
      RECT 0.935000  2.175000 1.320000 2.465000 ;
      RECT 1.150000  0.545000 1.320000 1.075000 ;
      RECT 1.150000  1.075000 1.900000 1.275000 ;
      RECT 1.150000  1.275000 1.320000 2.175000 ;
      RECT 1.515000  0.255000 1.740000 0.735000 ;
      RECT 1.515000  0.735000 2.240000 0.905000 ;
      RECT 1.515000  1.575000 2.240000 1.745000 ;
      RECT 1.515000  1.745000 1.740000 2.430000 ;
      RECT 1.910000  0.085000 2.240000 0.565000 ;
      RECT 1.910000  1.915000 2.270000 2.635000 ;
      RECT 2.070000  0.905000 2.240000 0.995000 ;
      RECT 2.070000  0.995000 2.360000 1.325000 ;
      RECT 2.070000  1.325000 2.240000 1.575000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__dlygate4sd1_1
MACRO sky130_fd_sc_hd__dlygate4sd2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlygate4sd2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.625000 1.615000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.570000 0.255000 3.135000 0.825000 ;
        RECT 2.570000 1.495000 3.135000 2.465000 ;
        RECT 2.675000 0.825000 3.135000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.255000 0.485000 0.715000 ;
      RECT 0.085000  0.715000 1.030000 0.885000 ;
      RECT 0.085000  1.785000 1.030000 2.005000 ;
      RECT 0.085000  2.005000 0.485000 2.465000 ;
      RECT 0.655000  0.085000 0.925000 0.545000 ;
      RECT 0.655000  2.175000 0.925000 2.635000 ;
      RECT 0.795000  0.885000 1.030000 0.995000 ;
      RECT 0.795000  0.995000 1.085000 1.325000 ;
      RECT 0.795000  1.325000 1.030000 1.785000 ;
      RECT 1.155000  0.255000 1.425000 0.585000 ;
      RECT 1.155000  2.135000 1.425000 2.465000 ;
      RECT 1.255000  0.585000 1.425000 1.055000 ;
      RECT 1.255000  1.055000 2.030000 1.615000 ;
      RECT 1.255000  1.615000 1.425000 2.135000 ;
      RECT 1.615000  0.255000 1.875000 0.715000 ;
      RECT 1.615000  0.715000 2.400000 0.885000 ;
      RECT 1.615000  1.785000 2.400000 2.005000 ;
      RECT 1.615000  2.005000 1.875000 2.465000 ;
      RECT 2.075000  0.085000 2.400000 0.545000 ;
      RECT 2.075000  2.175000 2.400000 2.635000 ;
      RECT 2.200000  0.885000 2.400000 0.995000 ;
      RECT 2.200000  0.995000 2.505000 1.325000 ;
      RECT 2.200000  1.325000 2.400000 1.785000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__dlygate4sd2_1
MACRO sky130_fd_sc_hd__dlygate4sd3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlygate4sd3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.775000 1.615000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.210000 0.255000 3.595000 0.825000 ;
        RECT 3.210000 1.495000 3.595000 2.465000 ;
        RECT 3.315000 0.825000 3.595000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.200000  0.255000 0.485000 0.715000 ;
      RECT 0.200000  0.715000 1.155000 0.885000 ;
      RECT 0.200000  1.785000 1.155000 2.005000 ;
      RECT 0.200000  2.005000 0.485000 2.465000 ;
      RECT 0.655000  0.085000 0.925000 0.545000 ;
      RECT 0.655000  2.175000 0.925000 2.635000 ;
      RECT 0.945000  0.885000 1.155000 1.785000 ;
      RECT 1.325000  0.255000 1.725000 1.055000 ;
      RECT 1.325000  1.055000 2.420000 1.615000 ;
      RECT 1.325000  1.615000 1.725000 2.465000 ;
      RECT 1.915000  0.255000 2.195000 0.715000 ;
      RECT 1.915000  0.715000 3.040000 0.885000 ;
      RECT 1.915000  1.785000 3.040000 2.005000 ;
      RECT 1.915000  2.005000 2.195000 2.465000 ;
      RECT 2.590000  0.885000 3.040000 0.995000 ;
      RECT 2.590000  0.995000 3.145000 1.325000 ;
      RECT 2.590000  1.325000 3.040000 1.785000 ;
      RECT 2.715000  0.085000 3.040000 0.545000 ;
      RECT 2.715000  2.175000 3.040000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__dlygate4sd3_1
MACRO sky130_fd_sc_hd__dlymetal6s2s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlymetal6s2s_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.570000 1.700000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.245000 0.255000 1.670000 0.825000 ;
        RECT 1.245000 1.495000 2.150000 1.675000 ;
        RECT 1.245000 1.675000 1.670000 2.465000 ;
        RECT 1.320000 0.825000 1.670000 0.995000 ;
        RECT 1.320000 0.995000 2.150000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.120000 -0.085000 0.290000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.255000 0.520000 0.655000 ;
      RECT 0.085000  0.655000 1.075000 0.825000 ;
      RECT 0.085000  1.870000 1.075000 2.040000 ;
      RECT 0.085000  2.040000 0.520000 2.465000 ;
      RECT 0.690000  0.085000 1.075000 0.485000 ;
      RECT 0.690000  2.210000 1.075000 2.635000 ;
      RECT 0.740000  0.825000 1.075000 0.995000 ;
      RECT 0.740000  0.995000 1.150000 1.325000 ;
      RECT 0.740000  1.325000 1.075000 1.870000 ;
      RECT 1.840000  1.845000 2.670000 2.040000 ;
      RECT 1.840000  2.040000 2.115000 2.465000 ;
      RECT 1.860000  0.255000 2.115000 0.655000 ;
      RECT 1.860000  0.655000 2.670000 0.825000 ;
      RECT 2.285000  0.085000 2.670000 0.485000 ;
      RECT 2.285000  2.210000 2.670000 2.635000 ;
      RECT 2.320000  0.825000 2.670000 0.995000 ;
      RECT 2.320000  0.995000 2.745000 1.325000 ;
      RECT 2.320000  1.325000 2.670000 1.845000 ;
      RECT 2.840000  0.255000 3.085000 0.825000 ;
      RECT 2.840000  1.495000 3.565000 1.675000 ;
      RECT 2.840000  1.675000 3.085000 2.465000 ;
      RECT 2.915000  0.825000 3.085000 0.995000 ;
      RECT 2.915000  0.995000 3.565000 1.495000 ;
      RECT 3.275000  0.255000 3.530000 0.655000 ;
      RECT 3.275000  0.655000 4.085000 0.825000 ;
      RECT 3.275000  1.845000 4.085000 2.040000 ;
      RECT 3.275000  2.040000 3.530000 2.465000 ;
      RECT 3.700000  0.085000 4.085000 0.485000 ;
      RECT 3.700000  2.210000 4.085000 2.635000 ;
      RECT 3.735000  0.825000 4.085000 0.995000 ;
      RECT 3.735000  0.995000 4.160000 1.325000 ;
      RECT 3.735000  1.325000 4.085000 1.845000 ;
      RECT 4.255000  0.255000 4.515000 0.825000 ;
      RECT 4.255000  1.495000 4.515000 2.465000 ;
      RECT 4.330000  0.825000 4.515000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__dlymetal6s2s_1
MACRO sky130_fd_sc_hd__dlymetal6s4s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlymetal6s4s_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.570000 1.700000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.660000 0.255000 3.105000 0.825000 ;
        RECT 2.660000 1.495000 3.565000 1.675000 ;
        RECT 2.660000 1.675000 3.105000 2.465000 ;
        RECT 2.735000 0.825000 3.105000 0.995000 ;
        RECT 2.735000 0.995000 3.565000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.120000 -0.085000 0.290000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.255000 0.520000 0.655000 ;
      RECT 0.085000  0.655000 1.075000 0.825000 ;
      RECT 0.085000  1.870000 1.075000 2.040000 ;
      RECT 0.085000  2.040000 0.520000 2.465000 ;
      RECT 0.690000  0.085000 1.075000 0.485000 ;
      RECT 0.690000  2.210000 1.075000 2.635000 ;
      RECT 0.740000  0.825000 1.075000 0.995000 ;
      RECT 0.740000  0.995000 1.150000 1.325000 ;
      RECT 0.740000  1.325000 1.075000 1.870000 ;
      RECT 1.245000  0.255000 1.515000 0.825000 ;
      RECT 1.245000  1.495000 1.970000 1.675000 ;
      RECT 1.245000  1.675000 1.515000 2.465000 ;
      RECT 1.320000  0.825000 1.515000 0.995000 ;
      RECT 1.320000  0.995000 1.970000 1.495000 ;
      RECT 1.685000  0.255000 1.935000 0.655000 ;
      RECT 1.685000  0.655000 2.490000 0.825000 ;
      RECT 1.685000  1.845000 2.490000 2.040000 ;
      RECT 1.685000  2.040000 1.935000 2.465000 ;
      RECT 2.105000  0.085000 2.490000 0.485000 ;
      RECT 2.105000  2.210000 2.490000 2.635000 ;
      RECT 2.140000  0.825000 2.490000 0.995000 ;
      RECT 2.140000  0.995000 2.565000 1.325000 ;
      RECT 2.140000  1.325000 2.490000 1.845000 ;
      RECT 3.275000  0.255000 3.530000 0.655000 ;
      RECT 3.275000  0.655000 4.085000 0.825000 ;
      RECT 3.275000  1.845000 4.085000 2.040000 ;
      RECT 3.275000  2.040000 3.530000 2.465000 ;
      RECT 3.700000  0.085000 4.085000 0.485000 ;
      RECT 3.700000  2.210000 4.085000 2.635000 ;
      RECT 3.735000  0.825000 4.085000 0.995000 ;
      RECT 3.735000  0.995000 4.160000 1.325000 ;
      RECT 3.735000  1.325000 4.085000 1.845000 ;
      RECT 4.255000  0.255000 4.515000 0.825000 ;
      RECT 4.255000  1.495000 4.515000 2.465000 ;
      RECT 4.330000  0.825000 4.515000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__dlymetal6s4s_1
MACRO sky130_fd_sc_hd__dlymetal6s6s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlymetal6s6s_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.575000 1.700000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.080000 0.255000 4.515000 0.825000 ;
        RECT 4.080000 1.495000 4.515000 2.465000 ;
        RECT 4.155000 0.825000 4.515000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.125000 -0.085000 0.295000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.255000 0.525000 0.655000 ;
      RECT 0.085000  0.655000 1.080000 0.825000 ;
      RECT 0.085000  1.870000 1.080000 2.040000 ;
      RECT 0.085000  2.040000 0.525000 2.465000 ;
      RECT 0.695000  0.085000 1.080000 0.485000 ;
      RECT 0.695000  2.210000 1.080000 2.635000 ;
      RECT 0.745000  0.825000 1.080000 0.995000 ;
      RECT 0.745000  0.995000 1.155000 1.325000 ;
      RECT 0.745000  1.325000 1.080000 1.870000 ;
      RECT 1.250000  0.255000 1.520000 0.825000 ;
      RECT 1.250000  1.495000 1.975000 1.675000 ;
      RECT 1.250000  1.675000 1.520000 2.465000 ;
      RECT 1.325000  0.825000 1.520000 0.995000 ;
      RECT 1.325000  0.995000 1.975000 1.495000 ;
      RECT 1.690000  0.255000 1.940000 0.655000 ;
      RECT 1.690000  0.655000 2.495000 0.825000 ;
      RECT 1.690000  1.845000 2.495000 2.040000 ;
      RECT 1.690000  2.040000 1.940000 2.465000 ;
      RECT 2.110000  0.085000 2.495000 0.485000 ;
      RECT 2.110000  2.210000 2.495000 2.635000 ;
      RECT 2.145000  0.825000 2.495000 0.995000 ;
      RECT 2.145000  0.995000 2.570000 1.325000 ;
      RECT 2.145000  1.325000 2.495000 1.845000 ;
      RECT 2.665000  0.255000 2.915000 0.825000 ;
      RECT 2.665000  1.495000 3.390000 1.675000 ;
      RECT 2.665000  1.675000 2.915000 2.465000 ;
      RECT 2.740000  0.825000 2.915000 0.995000 ;
      RECT 2.740000  0.995000 3.390000 1.495000 ;
      RECT 3.085000  0.255000 3.355000 0.655000 ;
      RECT 3.085000  0.655000 3.910000 0.825000 ;
      RECT 3.085000  1.845000 3.910000 2.040000 ;
      RECT 3.085000  2.040000 3.355000 2.465000 ;
      RECT 3.525000  0.085000 3.910000 0.485000 ;
      RECT 3.525000  2.210000 3.910000 2.635000 ;
      RECT 3.560000  0.825000 3.910000 0.995000 ;
      RECT 3.560000  0.995000 3.985000 1.325000 ;
      RECT 3.560000  1.325000 3.910000 1.845000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__dlymetal6s6s_1
MACRO sky130_fd_sc_hd__ebufn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.355000 1.615000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.309000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.910000 1.075000 1.240000 1.630000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.601000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.495000 3.595000 2.465000 ;
        RECT 3.125000 0.255000 3.595000 0.825000 ;
        RECT 3.255000 0.825000 3.595000 1.495000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.280000 0.345000 0.615000 ;
      RECT 0.085000  0.615000 1.185000 0.825000 ;
      RECT 0.085000  1.785000 0.740000 2.005000 ;
      RECT 0.085000  2.005000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.445000 ;
      RECT 0.515000  2.175000 0.845000 2.635000 ;
      RECT 0.525000  0.825000 0.740000 1.785000 ;
      RECT 1.015000  0.255000 2.025000 0.465000 ;
      RECT 1.015000  0.465000 1.185000 0.615000 ;
      RECT 1.015000  1.800000 1.805000 2.005000 ;
      RECT 1.015000  2.005000 1.270000 2.460000 ;
      RECT 1.355000  0.635000 1.685000 0.885000 ;
      RECT 1.410000  0.885000 1.685000 1.075000 ;
      RECT 1.410000  1.075000 2.535000 1.325000 ;
      RECT 1.410000  1.325000 1.805000 1.800000 ;
      RECT 1.440000  2.175000 1.805000 2.635000 ;
      RECT 1.855000  0.465000 2.025000 0.735000 ;
      RECT 1.855000  0.735000 2.955000 0.905000 ;
      RECT 2.195000  0.085000 2.955000 0.565000 ;
      RECT 2.705000  0.905000 2.955000 0.995000 ;
      RECT 2.705000  0.995000 3.085000 1.325000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__ebufn_1
MACRO sky130_fd_sc_hd__ebufn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.490000 0.765000 0.780000 1.675000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.441000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.765000 1.280000 1.275000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.905000 1.445000 4.055000 1.625000 ;
        RECT 1.905000 1.625000 3.625000 1.765000 ;
        RECT 3.295000 0.635000 4.055000 0.855000 ;
        RECT 3.295000 1.765000 3.625000 2.125000 ;
        RECT 3.825000 0.855000 4.055000 1.445000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.280000 0.345000 0.615000 ;
      RECT 0.085000  0.615000 0.320000 1.845000 ;
      RECT 0.085000  1.845000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.850000 0.595000 ;
      RECT 0.515000  1.845000 0.950000 2.635000 ;
      RECT 1.020000  0.255000 1.730000 0.595000 ;
      RECT 1.120000  1.445000 1.735000 1.765000 ;
      RECT 1.120000  1.765000 1.410000 2.465000 ;
      RECT 1.450000  0.595000 1.730000 1.025000 ;
      RECT 1.450000  1.025000 2.965000 1.275000 ;
      RECT 1.450000  1.275000 1.735000 1.445000 ;
      RECT 1.600000  1.935000 3.125000 2.105000 ;
      RECT 1.600000  2.105000 1.810000 2.465000 ;
      RECT 1.900000  0.255000 2.170000 0.655000 ;
      RECT 1.900000  0.655000 3.125000 0.855000 ;
      RECT 1.980000  2.275000 2.310000 2.635000 ;
      RECT 2.340000  0.085000 2.670000 0.485000 ;
      RECT 2.480000  2.105000 3.125000 2.295000 ;
      RECT 2.480000  2.295000 4.055000 2.465000 ;
      RECT 2.840000  0.275000 4.050000 0.465000 ;
      RECT 2.840000  0.465000 3.125000 0.655000 ;
      RECT 3.245000  1.025000 3.655000 1.275000 ;
      RECT 3.795000  1.795000 4.055000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.150000  1.105000 0.320000 1.275000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.380000  1.105000 3.550000 1.275000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
    LAYER met1 ;
      RECT 0.085000 1.075000 0.380000 1.120000 ;
      RECT 0.085000 1.120000 3.610000 1.260000 ;
      RECT 0.085000 1.260000 0.380000 1.305000 ;
      RECT 3.320000 1.075000 3.610000 1.120000 ;
      RECT 3.320000 1.260000 3.610000 1.305000 ;
  END
END sky130_fd_sc_hd__ebufn_2
MACRO sky130_fd_sc_hd__ebufn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.490000 0.765000 0.780000 1.675000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.811500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.765000 1.280000 1.425000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895000 1.445000 5.895000 1.725000 ;
        RECT 4.145000 0.615000 5.895000 0.855000 ;
        RECT 5.675000 0.855000 5.895000 1.445000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.280000 0.345000 0.665000 ;
      RECT 0.085000  0.665000 0.320000 1.765000 ;
      RECT 0.085000  1.765000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.930000 0.595000 ;
      RECT 0.515000  1.845000 0.930000 2.635000 ;
      RECT 1.100000  0.255000 1.725000 0.595000 ;
      RECT 1.100000  1.595000 1.725000 1.765000 ;
      RECT 1.100000  1.765000 1.355000 2.465000 ;
      RECT 1.450000  0.595000 1.725000 1.025000 ;
      RECT 1.450000  1.025000 3.810000 1.275000 ;
      RECT 1.450000  1.275000 1.725000 1.595000 ;
      RECT 1.565000  1.935000 5.895000 2.105000 ;
      RECT 1.565000  2.105000 1.810000 2.465000 ;
      RECT 1.895000  0.255000 2.175000 0.655000 ;
      RECT 1.895000  0.655000 3.975000 0.855000 ;
      RECT 1.895000  1.895000 5.895000 1.935000 ;
      RECT 1.980000  2.275000 2.310000 2.635000 ;
      RECT 2.345000  0.085000 2.675000 0.485000 ;
      RECT 2.480000  2.105000 2.650000 2.465000 ;
      RECT 2.820000  2.275000 3.150000 2.635000 ;
      RECT 2.845000  0.275000 3.015000 0.655000 ;
      RECT 3.185000  0.085000 3.515000 0.485000 ;
      RECT 3.320000  2.105000 5.895000 2.465000 ;
      RECT 3.685000  0.255000 5.735000 0.445000 ;
      RECT 3.685000  0.445000 3.975000 0.655000 ;
      RECT 3.980000  1.025000 5.505000 1.275000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.150000  1.105000 0.320000 1.275000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.310000  1.105000 4.480000 1.275000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 0.085000 1.075000 0.380000 1.120000 ;
      RECT 0.085000 1.120000 4.540000 1.260000 ;
      RECT 0.085000 1.260000 0.380000 1.305000 ;
      RECT 4.250000 1.075000 4.540000 1.120000 ;
      RECT 4.250000 1.260000 4.540000 1.305000 ;
  END
END sky130_fd_sc_hd__ebufn_4
MACRO sky130_fd_sc_hd__ebufn_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.430000 1.615000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.375500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.970000 0.620000 1.305000 0.995000 ;
        RECT 0.970000 0.995000 1.430000 1.325000 ;
        RECT 0.970000 1.325000 1.305000 1.695000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995000 1.445000 9.575000 1.725000 ;
        RECT 6.275000 0.615000 9.575000 0.855000 ;
        RECT 9.325000 0.855000 9.575000 1.445000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.085000  0.085000 0.445000 0.825000 ;
      RECT 0.085000  1.785000 0.445000 2.635000 ;
      RECT 0.600000  0.995000 0.800000 1.615000 ;
      RECT 0.615000  0.280000 0.800000 0.995000 ;
      RECT 0.615000  1.615000 0.800000 2.465000 ;
      RECT 0.970000  0.085000 1.305000 0.445000 ;
      RECT 0.970000  1.865000 1.305000 2.635000 ;
      RECT 1.475000  0.255000 1.985000 0.825000 ;
      RECT 1.475000  1.495000 1.825000 2.465000 ;
      RECT 1.600000  0.825000 1.985000 1.025000 ;
      RECT 1.600000  1.025000 5.925000 1.275000 ;
      RECT 1.600000  1.275000 1.825000 1.495000 ;
      RECT 1.995000  1.895000 9.575000 2.065000 ;
      RECT 1.995000  2.065000 2.245000 2.465000 ;
      RECT 2.155000  0.255000 2.485000 0.655000 ;
      RECT 2.155000  0.655000 6.105000 0.855000 ;
      RECT 2.415000  2.235000 2.745000 2.635000 ;
      RECT 2.655000  0.085000 2.985000 0.485000 ;
      RECT 2.915000  2.065000 3.085000 2.465000 ;
      RECT 3.155000  0.275000 3.325000 0.655000 ;
      RECT 3.255000  2.235000 3.585000 2.635000 ;
      RECT 3.495000  0.085000 3.825000 0.485000 ;
      RECT 3.755000  2.065000 3.925000 2.465000 ;
      RECT 3.995000  0.255000 4.165000 0.655000 ;
      RECT 4.095000  2.235000 4.425000 2.635000 ;
      RECT 4.335000  0.085000 4.665000 0.485000 ;
      RECT 4.595000  2.065000 4.765000 2.465000 ;
      RECT 4.835000  0.275000 5.005000 0.655000 ;
      RECT 4.935000  2.235000 5.265000 2.635000 ;
      RECT 5.175000  0.085000 5.505000 0.485000 ;
      RECT 5.435000  2.065000 9.575000 2.465000 ;
      RECT 5.675000  0.255000 9.575000 0.445000 ;
      RECT 5.675000  0.445000 6.105000 0.655000 ;
      RECT 6.175000  1.025000 9.155000 1.275000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  1.105000 0.775000 1.275000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.580000  1.105000 6.750000 1.275000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 0.545000 1.075000 0.835000 1.120000 ;
      RECT 0.545000 1.120000 6.810000 1.260000 ;
      RECT 0.545000 1.260000 0.835000 1.305000 ;
      RECT 6.520000 1.075000 6.810000 1.120000 ;
      RECT 6.520000 1.260000 6.810000 1.305000 ;
  END
END sky130_fd_sc_hd__ebufn_8
MACRO sky130_fd_sc_hd__edfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__edfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.765000 1.915000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 0.765000 2.565000 1.185000 ;
        RECT 2.110000 1.185000 2.325000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.225000 0.255000 11.555000 2.420000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.400000 1.065000 9.845000 1.410000 ;
        RECT 9.400000 1.410000 9.730000 2.465000 ;
        RECT 9.515000 0.255000 9.845000 1.065000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.150000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.845000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.355000  0.255000  1.785000 0.515000 ;
      RECT  1.355000  0.515000  1.525000 1.890000 ;
      RECT  1.355000  1.890000  1.785000 2.465000 ;
      RECT  2.235000  0.085000  2.565000 0.515000 ;
      RECT  2.235000  1.890000  2.565000 2.635000 ;
      RECT  2.495000  1.355000  3.085000 1.720000 ;
      RECT  2.755000  1.720000  3.085000 2.425000 ;
      RECT  2.780000  0.255000  3.005000 0.845000 ;
      RECT  2.780000  0.845000  3.635000 1.175000 ;
      RECT  2.780000  1.175000  3.085000 1.355000 ;
      RECT  3.185000  0.085000  3.515000 0.610000 ;
      RECT  3.265000  1.825000  3.460000 2.635000 ;
      RECT  3.805000  0.685000  3.975000 1.320000 ;
      RECT  3.805000  1.320000  4.175000 1.650000 ;
      RECT  4.125000  1.820000  4.515000 2.020000 ;
      RECT  4.125000  2.020000  4.455000 2.465000 ;
      RECT  4.145000  0.255000  4.415000 0.980000 ;
      RECT  4.145000  0.980000  4.515000 1.150000 ;
      RECT  4.345000  1.150000  4.515000 1.820000 ;
      RECT  4.795000  1.125000  4.980000 1.720000 ;
      RECT  4.815000  0.735000  5.320000 0.955000 ;
      RECT  4.915000  2.175000  5.955000 2.375000 ;
      RECT  5.005000  0.255000  5.680000 0.565000 ;
      RECT  5.150000  0.955000  5.320000 1.655000 ;
      RECT  5.150000  1.655000  5.615000 2.005000 ;
      RECT  5.510000  0.565000  5.680000 1.315000 ;
      RECT  5.510000  1.315000  6.360000 1.485000 ;
      RECT  5.785000  1.485000  6.360000 1.575000 ;
      RECT  5.785000  1.575000  5.955000 2.175000 ;
      RECT  5.870000  0.765000  6.935000 1.045000 ;
      RECT  5.870000  1.045000  7.445000 1.065000 ;
      RECT  5.870000  1.065000  6.070000 1.095000 ;
      RECT  5.945000  0.085000  6.340000 0.560000 ;
      RECT  6.125000  1.835000  6.360000 2.635000 ;
      RECT  6.190000  1.245000  6.360000 1.315000 ;
      RECT  6.530000  0.255000  6.935000 0.765000 ;
      RECT  6.530000  1.065000  7.445000 1.375000 ;
      RECT  6.530000  1.375000  6.860000 2.465000 ;
      RECT  7.070000  2.105000  7.360000 2.635000 ;
      RECT  7.165000  0.085000  7.440000 0.615000 ;
      RECT  7.790000  1.245000  7.980000 1.965000 ;
      RECT  7.925000  2.165000  8.890000 2.355000 ;
      RECT  8.005000  0.705000  8.470000 1.035000 ;
      RECT  8.025000  0.330000  8.890000 0.535000 ;
      RECT  8.150000  1.035000  8.470000 1.995000 ;
      RECT  8.640000  0.535000  8.890000 2.165000 ;
      RECT  9.060000  1.495000  9.230000 2.635000 ;
      RECT  9.095000  0.085000  9.345000 0.900000 ;
      RECT  9.900000  1.575000 10.130000 2.010000 ;
      RECT 10.015000  0.890000 10.640000 1.220000 ;
      RECT 10.300000  0.255000 10.640000 0.890000 ;
      RECT 10.300000  1.220000 10.640000 2.465000 ;
      RECT 10.810000  0.085000 11.055000 0.900000 ;
      RECT 10.810000  1.465000 11.055000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.635000  1.785000  0.805000 1.955000 ;
      RECT  1.015000  1.445000  1.185000 1.615000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.355000  0.425000  1.525000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.805000  0.765000  3.975000 0.935000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.185000  0.425000  4.355000 0.595000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.800000  1.445000  4.970000 1.615000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.210000  1.785000  5.380000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.800000  1.785000  7.970000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.220000  1.445000  8.390000 1.615000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.680000  1.785000  8.850000 1.955000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT  9.930000  1.785000 10.100000 1.955000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.390000  0.765000 10.560000 0.935000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
    LAYER met1 ;
      RECT  0.575000 1.755000  0.865000 1.800000 ;
      RECT  0.575000 1.800000  8.030000 1.940000 ;
      RECT  0.575000 1.940000  0.865000 1.985000 ;
      RECT  0.955000 1.415000  1.245000 1.460000 ;
      RECT  0.955000 1.460000  8.450000 1.600000 ;
      RECT  0.955000 1.600000  1.245000 1.645000 ;
      RECT  1.295000 0.395000  4.415000 0.580000 ;
      RECT  1.295000 0.580000  1.585000 0.625000 ;
      RECT  3.745000 0.735000  4.035000 0.780000 ;
      RECT  3.745000 0.780000 10.620000 0.920000 ;
      RECT  3.745000 0.920000  4.035000 0.965000 ;
      RECT  4.125000 0.580000  4.415000 0.625000 ;
      RECT  4.740000 1.415000  5.030000 1.460000 ;
      RECT  4.740000 1.600000  5.030000 1.645000 ;
      RECT  5.150000 1.755000  5.440000 1.800000 ;
      RECT  5.150000 1.940000  5.440000 1.985000 ;
      RECT  7.740000 1.755000  8.030000 1.800000 ;
      RECT  7.740000 1.940000  8.030000 1.985000 ;
      RECT  8.160000 1.415000  8.450000 1.460000 ;
      RECT  8.160000 1.600000  8.450000 1.645000 ;
      RECT  8.620000 1.755000  8.910000 1.800000 ;
      RECT  8.620000 1.800000 10.160000 1.940000 ;
      RECT  8.620000 1.940000  8.910000 1.985000 ;
      RECT  9.870000 1.755000 10.160000 1.800000 ;
      RECT  9.870000 1.940000 10.160000 1.985000 ;
      RECT 10.330000 0.735000 10.620000 0.780000 ;
      RECT 10.330000 0.920000 10.620000 0.965000 ;
  END
END sky130_fd_sc_hd__edfxbp_1
MACRO sky130_fd_sc_hd__edfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__edfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.765000 1.915000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 0.765000 2.565000 1.185000 ;
        RECT 2.110000 1.185000 2.325000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.465000 0.305000 10.795000 2.420000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.845000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.355000  0.255000  1.785000 0.515000 ;
      RECT  1.355000  0.515000  1.525000 1.890000 ;
      RECT  1.355000  1.890000  1.785000 2.465000 ;
      RECT  2.235000  0.085000  2.565000 0.515000 ;
      RECT  2.235000  1.890000  2.565000 2.635000 ;
      RECT  2.495000  1.355000  3.085000 1.720000 ;
      RECT  2.755000  1.720000  3.085000 2.425000 ;
      RECT  2.780000  0.255000  3.005000 0.845000 ;
      RECT  2.780000  0.845000  3.635000 1.175000 ;
      RECT  2.780000  1.175000  3.085000 1.355000 ;
      RECT  3.185000  0.085000  3.515000 0.610000 ;
      RECT  3.265000  1.825000  3.460000 2.635000 ;
      RECT  3.805000  0.685000  3.975000 1.320000 ;
      RECT  3.805000  1.320000  4.175000 1.650000 ;
      RECT  4.125000  1.820000  4.515000 2.020000 ;
      RECT  4.125000  2.020000  4.455000 2.465000 ;
      RECT  4.145000  0.255000  4.415000 0.980000 ;
      RECT  4.145000  0.980000  4.515000 1.150000 ;
      RECT  4.345000  1.150000  4.515000 1.820000 ;
      RECT  4.795000  1.125000  4.980000 1.720000 ;
      RECT  4.815000  0.735000  5.320000 0.955000 ;
      RECT  4.915000  2.175000  5.955000 2.375000 ;
      RECT  5.005000  0.255000  5.680000 0.565000 ;
      RECT  5.150000  0.955000  5.320000 1.655000 ;
      RECT  5.150000  1.655000  5.615000 2.005000 ;
      RECT  5.510000  0.565000  5.680000 1.315000 ;
      RECT  5.510000  1.315000  6.360000 1.485000 ;
      RECT  5.785000  1.485000  6.360000 1.575000 ;
      RECT  5.785000  1.575000  5.955000 2.175000 ;
      RECT  5.870000  0.765000  6.935000 1.045000 ;
      RECT  5.870000  1.045000  7.445000 1.065000 ;
      RECT  5.870000  1.065000  6.070000 1.095000 ;
      RECT  5.945000  0.085000  6.340000 0.560000 ;
      RECT  6.125000  1.835000  6.360000 2.635000 ;
      RECT  6.190000  1.245000  6.360000 1.315000 ;
      RECT  6.530000  0.255000  6.935000 0.765000 ;
      RECT  6.530000  1.065000  7.445000 1.375000 ;
      RECT  6.530000  1.375000  6.860000 2.465000 ;
      RECT  7.070000  2.105000  7.360000 2.635000 ;
      RECT  7.165000  0.085000  7.440000 0.615000 ;
      RECT  7.790000  1.245000  7.980000 1.965000 ;
      RECT  7.925000  2.165000  8.810000 2.355000 ;
      RECT  8.005000  0.705000  8.470000 1.035000 ;
      RECT  8.025000  0.330000  8.810000 0.535000 ;
      RECT  8.150000  1.035000  8.470000 1.995000 ;
      RECT  8.640000  0.535000  8.810000 0.995000 ;
      RECT  8.640000  0.995000  9.510000 1.325000 ;
      RECT  8.640000  1.325000  8.810000 2.165000 ;
      RECT  8.980000  1.530000  9.880000 1.905000 ;
      RECT  8.980000  2.135000  9.240000 2.635000 ;
      RECT  9.050000  0.085000  9.365000 0.615000 ;
      RECT  9.540000  1.905000  9.880000 2.465000 ;
      RECT  9.550000  0.300000  9.880000 0.825000 ;
      RECT  9.690000  0.825000  9.880000 1.530000 ;
      RECT 10.050000  0.085000 10.295000 0.900000 ;
      RECT 10.050000  1.465000 10.295000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.635000  1.785000  0.805000 1.955000 ;
      RECT  1.015000  1.445000  1.185000 1.615000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.355000  0.425000  1.525000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.805000  0.765000  3.975000 0.935000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.185000  0.425000  4.355000 0.595000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.800000  1.445000  4.970000 1.615000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.210000  1.785000  5.380000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.800000  1.785000  7.970000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.220000  1.445000  8.390000 1.615000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.700000  0.765000  9.870000 0.935000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 0.575000 1.755000 0.865000 1.800000 ;
      RECT 0.575000 1.800000 8.030000 1.940000 ;
      RECT 0.575000 1.940000 0.865000 1.985000 ;
      RECT 0.955000 1.415000 1.245000 1.460000 ;
      RECT 0.955000 1.460000 8.450000 1.600000 ;
      RECT 0.955000 1.600000 1.245000 1.645000 ;
      RECT 1.295000 0.395000 4.415000 0.580000 ;
      RECT 1.295000 0.580000 1.585000 0.625000 ;
      RECT 3.745000 0.735000 4.035000 0.780000 ;
      RECT 3.745000 0.780000 9.930000 0.920000 ;
      RECT 3.745000 0.920000 4.035000 0.965000 ;
      RECT 4.125000 0.580000 4.415000 0.625000 ;
      RECT 4.740000 1.415000 5.030000 1.460000 ;
      RECT 4.740000 1.600000 5.030000 1.645000 ;
      RECT 5.150000 1.755000 5.440000 1.800000 ;
      RECT 5.150000 1.940000 5.440000 1.985000 ;
      RECT 7.740000 1.755000 8.030000 1.800000 ;
      RECT 7.740000 1.940000 8.030000 1.985000 ;
      RECT 8.160000 1.415000 8.450000 1.460000 ;
      RECT 8.160000 1.600000 8.450000 1.645000 ;
      RECT 9.640000 0.735000 9.930000 0.780000 ;
      RECT 9.640000 0.920000 9.930000 0.965000 ;
  END
END sky130_fd_sc_hd__edfxtp_1
MACRO sky130_fd_sc_hd__einvn_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 0.765000 1.755000 1.955000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.650000 1.725000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.275600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.160000 0.255000 1.755000 0.595000 ;
        RECT 1.160000 0.595000 1.330000 2.125000 ;
        RECT 1.160000 2.125000 1.755000 2.465000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.085000  0.255000 0.360000 0.655000 ;
      RECT 0.085000  0.655000 0.990000 0.825000 ;
      RECT 0.085000  1.895000 0.990000 2.065000 ;
      RECT 0.085000  2.065000 0.400000 2.465000 ;
      RECT 0.530000  0.085000 0.990000 0.485000 ;
      RECT 0.570000  2.235000 0.990000 2.635000 ;
      RECT 0.820000  0.825000 0.990000 1.895000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__einvn_0
MACRO sky130_fd_sc_hd__einvn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.970000 0.765000 2.215000 1.615000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.309000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.510000 1.725000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.040000 1.785000 2.215000 2.465000 ;
        RECT 1.620000 0.255000 2.215000 0.595000 ;
        RECT 1.620000 0.595000 1.800000 1.785000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.085000  0.255000 0.370000 0.615000 ;
      RECT 0.085000  0.615000 1.450000 0.785000 ;
      RECT 0.085000  1.895000 0.870000 2.065000 ;
      RECT 0.085000  2.065000 0.370000 2.465000 ;
      RECT 0.540000  0.085000 1.440000 0.445000 ;
      RECT 0.540000  2.235000 0.870000 2.635000 ;
      RECT 0.685000  0.785000 1.450000 1.615000 ;
      RECT 0.685000  1.615000 0.870000 1.895000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__einvn_1
MACRO sky130_fd_sc_hd__einvn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 1.075000 3.135000 1.275000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.441000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.325000 1.385000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.694800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 1.445000 3.135000 1.695000 ;
        RECT 2.365000 0.595000 2.695000 0.845000 ;
        RECT 2.365000 0.845000 2.615000 1.445000 ;
        RECT 2.785000 1.695000 3.135000 2.465000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.840000 0.825000 ;
      RECT 0.085000  1.555000 0.895000 1.725000 ;
      RECT 0.085000  1.725000 0.345000 2.465000 ;
      RECT 0.495000  0.825000 0.840000 0.995000 ;
      RECT 0.495000  0.995000 2.035000 1.275000 ;
      RECT 0.495000  1.275000 0.895000 1.555000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 0.515000  1.895000 0.895000 2.635000 ;
      RECT 1.015000  0.255000 1.280000 0.655000 ;
      RECT 1.015000  0.655000 2.195000 0.825000 ;
      RECT 1.070000  1.445000 1.775000 1.865000 ;
      RECT 1.070000  1.865000 2.615000 2.085000 ;
      RECT 1.070000  2.085000 1.240000 2.465000 ;
      RECT 1.410000  2.255000 2.275000 2.635000 ;
      RECT 1.450000  0.085000 1.780000 0.485000 ;
      RECT 1.950000  0.255000 3.135000 0.425000 ;
      RECT 1.950000  0.425000 2.195000 0.655000 ;
      RECT 2.445000  2.085000 2.615000 2.465000 ;
      RECT 2.865000  0.425000 3.135000 0.775000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__einvn_2
MACRO sky130_fd_sc_hd__einvn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.530000 0.620000 4.975000 1.325000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.811500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.345000 1.325000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.190000 0.620000 4.360000 1.480000 ;
        RECT 3.190000 1.480000 3.520000 2.075000 ;
        RECT 4.030000 1.480000 4.360000 2.075000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.845000 0.825000 ;
      RECT 0.085000  1.495000 0.845000 1.665000 ;
      RECT 0.085000  1.665000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 0.515000  0.825000 0.845000 0.995000 ;
      RECT 0.515000  0.995000 3.020000 1.325000 ;
      RECT 0.515000  1.325000 0.845000 1.495000 ;
      RECT 0.515000  1.835000 0.845000 2.635000 ;
      RECT 1.015000  0.255000 1.285000 0.655000 ;
      RECT 1.015000  0.655000 2.995000 0.825000 ;
      RECT 1.015000  1.495000 3.020000 1.665000 ;
      RECT 1.015000  1.665000 1.240000 2.465000 ;
      RECT 1.410000  1.835000 1.740000 2.635000 ;
      RECT 1.455000  0.085000 1.785000 0.485000 ;
      RECT 1.910000  1.665000 2.080000 2.465000 ;
      RECT 1.955000  0.255000 2.125000 0.655000 ;
      RECT 2.250000  1.835000 2.640000 2.635000 ;
      RECT 2.295000  0.085000 2.625000 0.485000 ;
      RECT 2.810000  1.665000 3.020000 2.295000 ;
      RECT 2.810000  2.295000 4.975000 2.465000 ;
      RECT 2.825000  0.255000 4.975000 0.450000 ;
      RECT 2.825000  0.450000 2.995000 0.655000 ;
      RECT 3.690000  1.650000 3.860000 2.295000 ;
      RECT 4.530000  1.650000 4.975000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__einvn_4
MACRO sky130_fd_sc_hd__einvn_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.645000 0.995000 7.800000 1.285000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.375500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.345000 1.325000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.870000 0.620000 8.195000 0.825000 ;
        RECT 4.870000 1.455000 8.195000 1.625000 ;
        RECT 4.870000 1.625000 5.200000 2.125000 ;
        RECT 5.710000 1.625000 6.040000 2.125000 ;
        RECT 6.550000 1.625000 6.880000 2.125000 ;
        RECT 7.390000 1.625000 7.720000 2.125000 ;
        RECT 7.970000 0.825000 8.195000 1.455000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.090000  0.255000 0.345000 0.655000 ;
      RECT 0.090000  0.655000 0.845000 0.825000 ;
      RECT 0.090000  1.495000 0.845000 1.665000 ;
      RECT 0.090000  1.665000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 0.515000  0.825000 0.845000 0.995000 ;
      RECT 0.515000  0.995000 4.475000 1.325000 ;
      RECT 0.515000  1.325000 0.845000 1.495000 ;
      RECT 0.515000  1.835000 0.845000 2.635000 ;
      RECT 1.015000  0.255000 1.285000 0.655000 ;
      RECT 1.015000  0.655000 4.700000 0.825000 ;
      RECT 1.015000  1.495000 4.700000 1.665000 ;
      RECT 1.015000  1.665000 1.240000 2.465000 ;
      RECT 1.410000  1.835000 1.740000 2.635000 ;
      RECT 1.455000  0.085000 1.785000 0.485000 ;
      RECT 1.910000  1.665000 2.080000 2.465000 ;
      RECT 1.955000  0.255000 2.125000 0.655000 ;
      RECT 2.250000  1.835000 2.580000 2.635000 ;
      RECT 2.295000  0.085000 2.625000 0.485000 ;
      RECT 2.750000  1.665000 2.920000 2.465000 ;
      RECT 2.795000  0.255000 2.965000 0.655000 ;
      RECT 3.090000  1.835000 3.420000 2.635000 ;
      RECT 3.135000  0.085000 3.465000 0.485000 ;
      RECT 3.590000  1.665000 3.760000 2.465000 ;
      RECT 3.635000  0.255000 3.805000 0.655000 ;
      RECT 3.930000  1.835000 4.280000 2.635000 ;
      RECT 3.975000  0.085000 4.315000 0.485000 ;
      RECT 4.450000  1.665000 4.700000 2.295000 ;
      RECT 4.450000  2.295000 8.195000 2.465000 ;
      RECT 4.485000  0.255000 8.195000 0.450000 ;
      RECT 4.485000  0.450000 4.700000 0.655000 ;
      RECT 5.370000  1.795000 5.540000 2.295000 ;
      RECT 6.210000  1.795000 6.380000 2.295000 ;
      RECT 7.050000  1.795000 7.220000 2.295000 ;
      RECT 7.890000  1.795000 8.195000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
END sky130_fd_sc_hd__einvn_8
MACRO sky130_fd_sc_hd__einvp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 0.975000 2.215000 1.955000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.223500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.545000 1.725000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.620000 0.255000 2.215000 0.805000 ;
        RECT 1.620000 0.805000 1.795000 2.125000 ;
        RECT 1.620000 2.125000 2.215000 2.465000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 1.450000 0.825000 ;
      RECT 0.085000  1.895000 1.450000 2.065000 ;
      RECT 0.085000  2.065000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 1.450000 0.485000 ;
      RECT 0.515000  2.235000 1.450000 2.635000 ;
      RECT 0.715000  0.825000 1.450000 1.895000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__einvp_1
MACRO sky130_fd_sc_hd__einvp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.850000 0.765000 3.135000 1.615000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.354000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.330000 1.615000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.350000 0.595000 2.680000 2.125000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.875000 0.825000 ;
      RECT 0.085000  1.785000 0.875000 1.955000 ;
      RECT 0.085000  1.955000 0.345000 2.465000 ;
      RECT 0.500000  0.825000 0.875000 0.995000 ;
      RECT 0.500000  0.995000 2.180000 1.325000 ;
      RECT 0.500000  1.325000 0.875000 1.785000 ;
      RECT 0.515000  0.085000 0.875000 0.485000 ;
      RECT 0.515000  2.125000 0.875000 2.635000 ;
      RECT 1.045000  0.255000 1.240000 0.655000 ;
      RECT 1.045000  0.655000 2.180000 0.825000 ;
      RECT 1.045000  1.555000 2.155000 1.725000 ;
      RECT 1.045000  1.725000 1.285000 2.465000 ;
      RECT 1.410000  0.085000 1.770000 0.485000 ;
      RECT 1.455000  1.895000 1.785000 2.635000 ;
      RECT 1.940000  0.255000 3.135000 0.425000 ;
      RECT 1.940000  0.425000 2.180000 0.655000 ;
      RECT 1.985000  1.725000 2.155000 2.295000 ;
      RECT 1.985000  2.295000 3.135000 2.465000 ;
      RECT 2.850000  0.425000 3.135000 0.595000 ;
      RECT 2.850000  1.785000 3.135000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__einvp_2
MACRO sky130_fd_sc_hd__einvp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.740000 1.020000 4.975000 1.275000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.637500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.330000 1.615000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.190000 0.635000 4.975000 0.850000 ;
        RECT 3.190000 0.850000 3.570000 1.445000 ;
        RECT 3.190000 1.445000 4.360000 1.615000 ;
        RECT 3.190000 1.615000 3.520000 2.125000 ;
        RECT 4.030000 1.615000 4.360000 2.125000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.695000 0.825000 ;
      RECT 0.085000  1.785000 0.875000 1.955000 ;
      RECT 0.085000  1.955000 0.345000 2.465000 ;
      RECT 0.500000  0.825000 0.695000 0.995000 ;
      RECT 0.500000  0.995000 3.020000 1.325000 ;
      RECT 0.500000  1.325000 0.875000 1.785000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 0.515000  2.125000 0.875000 2.635000 ;
      RECT 1.035000  0.255000 1.205000 0.655000 ;
      RECT 1.035000  0.655000 3.020000 0.825000 ;
      RECT 1.075000  1.555000 2.995000 1.725000 ;
      RECT 1.075000  1.725000 1.285000 2.465000 ;
      RECT 1.375000  0.085000 1.705000 0.485000 ;
      RECT 1.455000  1.895000 1.785000 2.635000 ;
      RECT 1.875000  0.255000 2.045000 0.655000 ;
      RECT 1.955000  1.725000 2.125000 2.465000 ;
      RECT 2.215000  0.085000 2.555000 0.485000 ;
      RECT 2.295000  1.895000 2.655000 2.635000 ;
      RECT 2.735000  0.255000 4.975000 0.465000 ;
      RECT 2.735000  0.465000 3.020000 0.655000 ;
      RECT 2.825000  1.725000 2.995000 2.295000 ;
      RECT 2.825000  2.295000 4.975000 2.465000 ;
      RECT 3.690000  1.785000 3.860000 2.295000 ;
      RECT 4.530000  1.445000 4.975000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__einvp_4
MACRO sky130_fd_sc_hd__einvp_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.420000 1.020000 8.195000 1.275000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  1.027500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.330000 1.615000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.870000 0.635000 8.195000 0.850000 ;
        RECT 4.870000 0.850000 5.250000 1.445000 ;
        RECT 4.870000 1.445000 7.720000 1.615000 ;
        RECT 4.870000 1.615000 5.200000 2.125000 ;
        RECT 5.710000 1.615000 6.040000 2.125000 ;
        RECT 6.550000 1.615000 6.880000 2.125000 ;
        RECT 7.390000 1.615000 7.720000 2.125000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.695000 0.825000 ;
      RECT 0.085000  1.785000 0.875000 1.955000 ;
      RECT 0.085000  1.955000 0.345000 2.465000 ;
      RECT 0.500000  0.825000 0.695000 0.995000 ;
      RECT 0.500000  0.995000 4.700000 1.325000 ;
      RECT 0.500000  1.325000 0.875000 1.785000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 0.515000  2.125000 0.875000 2.635000 ;
      RECT 1.035000  0.255000 1.205000 0.655000 ;
      RECT 1.035000  0.655000 4.700000 0.825000 ;
      RECT 1.075000  1.555000 4.700000 1.725000 ;
      RECT 1.075000  1.725000 1.285000 2.465000 ;
      RECT 1.375000  0.085000 1.705000 0.485000 ;
      RECT 1.455000  1.895000 1.785000 2.635000 ;
      RECT 1.875000  0.255000 2.045000 0.655000 ;
      RECT 1.955000  1.725000 2.125000 2.465000 ;
      RECT 2.215000  0.085000 2.545000 0.485000 ;
      RECT 2.295000  1.895000 2.625000 2.635000 ;
      RECT 2.715000  0.255000 2.885000 0.655000 ;
      RECT 2.795000  1.725000 2.965000 2.465000 ;
      RECT 3.055000  0.085000 3.385000 0.485000 ;
      RECT 3.135000  1.895000 3.465000 2.635000 ;
      RECT 3.555000  0.255000 3.725000 0.655000 ;
      RECT 3.635000  1.725000 3.805000 2.465000 ;
      RECT 3.895000  0.085000 4.235000 0.485000 ;
      RECT 3.975000  1.895000 4.305000 2.635000 ;
      RECT 4.405000  0.255000 8.195000 0.465000 ;
      RECT 4.405000  0.465000 4.700000 0.655000 ;
      RECT 4.475000  1.725000 4.700000 2.295000 ;
      RECT 4.475000  2.295000 8.195000 2.465000 ;
      RECT 5.370000  1.785000 5.540000 2.295000 ;
      RECT 6.210000  1.785000 6.380000 2.295000 ;
      RECT 7.050000  1.785000 7.220000 2.295000 ;
      RECT 7.890000  1.445000 8.195000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
END sky130_fd_sc_hd__einvp_8
MACRO sky130_fd_sc_hd__fa_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fa_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.910000 0.995000 1.240000 1.275000 ;
        RECT 0.910000 1.275000 1.080000 1.325000 ;
      LAYER mcon ;
        RECT 1.070000 1.105000 1.240000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.230000 1.030000 2.620000 1.360000 ;
      LAYER mcon ;
        RECT 2.450000 1.105000 2.620000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.250000 0.955000 4.625000 1.275000 ;
      LAYER mcon ;
        RECT 4.310000 1.105000 4.480000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.885000 1.035000 6.325000 1.275000 ;
      LAYER mcon ;
        RECT 6.150000 1.105000 6.320000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.010000 1.075000 1.300000 1.120000 ;
        RECT 1.010000 1.120000 6.380000 1.260000 ;
        RECT 1.010000 1.260000 1.300000 1.305000 ;
        RECT 2.390000 1.075000 2.680000 1.120000 ;
        RECT 2.390000 1.260000 2.680000 1.305000 ;
        RECT 4.250000 1.075000 4.540000 1.120000 ;
        RECT 4.250000 1.260000 4.540000 1.305000 ;
        RECT 6.090000 1.075000 6.380000 1.120000 ;
        RECT 6.090000 1.260000 6.380000 1.305000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.300000 1.445000 1.700000 1.880000 ;
      LAYER mcon ;
        RECT 1.530000 1.445000 1.700000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.200000 1.435000 3.560000 1.765000 ;
      LAYER mcon ;
        RECT 3.390000 1.445000 3.560000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.635000 1.445000 6.055000 1.765000 ;
      LAYER mcon ;
        RECT 5.690000 1.445000 5.860000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.470000 1.415000 1.760000 1.460000 ;
        RECT 1.470000 1.460000 5.920000 1.600000 ;
        RECT 1.470000 1.600000 1.760000 1.645000 ;
        RECT 3.330000 1.415000 3.620000 1.460000 ;
        RECT 3.330000 1.600000 3.620000 1.645000 ;
        RECT 5.630000 1.415000 5.920000 1.460000 ;
        RECT 5.630000 1.600000 5.920000 1.645000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.670000 1.105000 2.040000 1.275000 ;
        RECT 1.870000 1.275000 2.040000 1.595000 ;
        RECT 1.870000 1.595000 2.960000 1.765000 ;
        RECT 2.790000 0.965000 3.955000 1.250000 ;
        RECT 2.790000 1.250000 2.960000 1.595000 ;
        RECT 3.785000 1.250000 3.955000 1.515000 ;
        RECT 3.785000 1.515000 5.405000 1.685000 ;
        RECT 5.155000 1.685000 5.405000 1.955000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.345000 0.830000 ;
        RECT 0.085000 0.830000 0.260000 1.485000 ;
        RECT 0.085000 1.485000 0.345000 2.465000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.840000 0.255000 7.240000 0.810000 ;
        RECT 6.840000 1.485000 7.240000 2.465000 ;
        RECT 6.910000 0.810000 7.240000 1.485000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.430000  0.995000 0.685000 1.325000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  0.635000 1.710000 0.805000 ;
      RECT 0.515000  0.805000 0.685000 0.995000 ;
      RECT 0.515000  1.325000 0.685000 1.625000 ;
      RECT 0.515000  1.625000 1.105000 1.945000 ;
      RECT 0.515000  2.150000 0.765000 2.635000 ;
      RECT 0.935000  1.945000 1.105000 2.065000 ;
      RECT 0.935000  2.065000 1.710000 2.465000 ;
      RECT 1.110000  0.255000 1.710000 0.635000 ;
      RECT 1.470000  0.805000 1.710000 0.935000 ;
      RECT 1.960000  0.255000 2.130000 0.615000 ;
      RECT 1.960000  0.615000 2.970000 0.785000 ;
      RECT 1.960000  1.935000 3.035000 2.105000 ;
      RECT 1.960000  2.105000 2.130000 2.465000 ;
      RECT 2.300000  0.085000 2.630000 0.445000 ;
      RECT 2.300000  2.275000 2.630000 2.635000 ;
      RECT 2.800000  0.255000 2.970000 0.615000 ;
      RECT 2.800000  2.105000 3.035000 2.465000 ;
      RECT 3.240000  0.085000 3.570000 0.490000 ;
      RECT 3.240000  2.255000 3.570000 2.635000 ;
      RECT 3.740000  0.255000 3.910000 0.615000 ;
      RECT 3.740000  0.615000 4.750000 0.785000 ;
      RECT 3.740000  1.935000 4.750000 2.105000 ;
      RECT 3.740000  2.105000 3.910000 2.465000 ;
      RECT 4.080000  0.085000 4.410000 0.445000 ;
      RECT 4.080000  2.275000 4.410000 2.635000 ;
      RECT 4.580000  0.255000 4.750000 0.615000 ;
      RECT 4.580000  2.105000 4.750000 2.465000 ;
      RECT 4.795000  0.955000 5.460000 1.125000 ;
      RECT 4.965000  0.765000 5.460000 0.955000 ;
      RECT 5.085000  0.255000 6.095000 0.505000 ;
      RECT 5.085000  0.505000 5.255000 0.595000 ;
      RECT 5.085000  2.125000 6.170000 2.465000 ;
      RECT 5.925000  0.505000 6.095000 0.615000 ;
      RECT 5.925000  0.615000 6.665000 0.785000 ;
      RECT 6.000000  1.935000 6.665000 2.105000 ;
      RECT 6.000000  2.105000 6.170000 2.125000 ;
      RECT 6.265000  0.085000 6.595000 0.445000 ;
      RECT 6.340000  2.275000 6.670000 2.635000 ;
      RECT 6.495000  0.785000 6.665000 0.995000 ;
      RECT 6.495000  0.995000 6.740000 1.325000 ;
      RECT 6.495000  1.325000 6.665000 1.935000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.530000  0.765000 1.700000 0.935000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.230000  0.765000 5.400000 0.935000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
    LAYER met1 ;
      RECT 1.470000 0.735000 1.760000 0.780000 ;
      RECT 1.470000 0.780000 5.460000 0.920000 ;
      RECT 1.470000 0.920000 1.760000 0.965000 ;
      RECT 5.170000 0.735000 5.460000 0.780000 ;
      RECT 5.170000 0.920000 5.460000 0.965000 ;
  END
END sky130_fd_sc_hd__fa_1
MACRO sky130_fd_sc_hd__fa_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fa_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.631500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.245000 0.995000 1.755000 1.275000 ;
        RECT 1.245000 1.275000 1.505000 1.325000 ;
      LAYER mcon ;
        RECT 1.525000 1.105000 1.695000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.685000 1.030000 3.075000 1.360000 ;
      LAYER mcon ;
        RECT 2.905000 1.105000 3.075000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.720000 0.955000 5.080000 1.275000 ;
      LAYER mcon ;
        RECT 4.765000 1.105000 4.935000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.105000 0.995000 6.960000 1.275000 ;
      LAYER mcon ;
        RECT 6.145000 1.105000 6.315000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465000 1.075000 1.755000 1.120000 ;
        RECT 1.465000 1.120000 6.375000 1.260000 ;
        RECT 1.465000 1.260000 1.755000 1.305000 ;
        RECT 2.845000 1.075000 3.135000 1.120000 ;
        RECT 2.845000 1.260000 3.135000 1.305000 ;
        RECT 4.705000 1.075000 4.995000 1.120000 ;
        RECT 4.705000 1.260000 4.995000 1.305000 ;
        RECT 6.085000 1.075000 6.375000 1.120000 ;
        RECT 6.085000 1.260000 6.375000 1.305000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.631500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.645000 1.445000 2.155000 1.690000 ;
      LAYER mcon ;
        RECT 1.985000 1.445000 2.155000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.655000 1.435000 4.070000 1.745000 ;
      LAYER mcon ;
        RECT 3.845000 1.445000 4.015000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.150000 1.445000 6.835000 1.735000 ;
      LAYER mcon ;
        RECT 6.605000 1.445000 6.775000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.925000 1.415000 2.215000 1.460000 ;
        RECT 1.925000 1.460000 6.835000 1.600000 ;
        RECT 1.925000 1.600000 2.215000 1.645000 ;
        RECT 3.785000 1.415000 4.075000 1.460000 ;
        RECT 3.785000 1.600000 4.075000 1.645000 ;
        RECT 6.545000 1.415000 6.835000 1.460000 ;
        RECT 6.545000 1.600000 6.835000 1.645000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.475500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.125000 1.105000 2.495000 1.275000 ;
        RECT 2.325000 1.275000 2.495000 1.570000 ;
        RECT 2.325000 1.570000 3.415000 1.740000 ;
        RECT 3.245000 0.965000 4.465000 1.250000 ;
        RECT 3.245000 1.250000 3.415000 1.570000 ;
        RECT 4.295000 1.250000 4.465000 1.435000 ;
        RECT 4.295000 1.435000 4.655000 1.515000 ;
        RECT 4.295000 1.515000 5.920000 1.685000 ;
        RECT 5.670000 1.355000 5.920000 1.515000 ;
        RECT 5.670000 1.685000 5.920000 1.955000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.735000 0.690000 0.905000 ;
        RECT 0.085000 0.905000 0.370000 1.415000 ;
        RECT 0.085000 1.415000 0.735000 1.585000 ;
        RECT 0.520000 0.315000 0.850000 0.485000 ;
        RECT 0.520000 0.485000 0.690000 0.735000 ;
        RECT 0.565000 1.585000 0.735000 1.780000 ;
        RECT 0.565000 1.780000 0.810000 1.950000 ;
        RECT 0.600000 1.950000 0.810000 2.465000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.523500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.395000 0.255000 7.725000 0.485000 ;
        RECT 7.395000 1.795000 7.645000 1.965000 ;
        RECT 7.395000 1.965000 7.565000 2.465000 ;
        RECT 7.475000 0.485000 7.725000 0.735000 ;
        RECT 7.475000 0.735000 8.195000 0.905000 ;
        RECT 7.475000 1.415000 8.195000 1.585000 ;
        RECT 7.475000 1.585000 7.645000 1.795000 ;
        RECT 7.970000 0.905000 8.195000 1.415000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.180000  0.085000 0.350000 0.565000 ;
      RECT 0.180000  1.795000 0.350000 2.635000 ;
      RECT 0.540000  1.075000 1.075000 1.245000 ;
      RECT 0.905000  0.655000 2.165000 0.825000 ;
      RECT 0.905000  0.825000 1.075000 1.075000 ;
      RECT 0.905000  1.245000 1.075000 1.430000 ;
      RECT 0.905000  1.430000 1.110000 1.495000 ;
      RECT 0.905000  1.495000 1.475000 1.600000 ;
      RECT 0.940000  1.600000 1.475000 1.665000 ;
      RECT 0.980000  2.275000 1.310000 2.635000 ;
      RECT 1.020000  0.085000 1.350000 0.465000 ;
      RECT 1.305000  1.665000 1.475000 1.910000 ;
      RECT 1.305000  1.910000 2.245000 2.080000 ;
      RECT 1.535000  0.255000 2.165000 0.655000 ;
      RECT 1.900000  2.080000 2.245000 2.465000 ;
      RECT 1.925000  0.825000 2.165000 0.935000 ;
      RECT 2.415000  0.255000 2.585000 0.615000 ;
      RECT 2.415000  0.615000 3.425000 0.785000 ;
      RECT 2.415000  1.935000 3.490000 2.105000 ;
      RECT 2.415000  2.105000 2.585000 2.465000 ;
      RECT 2.755000  0.085000 3.085000 0.445000 ;
      RECT 2.755000  2.275000 3.085000 2.635000 ;
      RECT 3.255000  0.255000 3.425000 0.615000 ;
      RECT 3.255000  2.105000 3.490000 2.465000 ;
      RECT 3.695000  0.085000 4.025000 0.490000 ;
      RECT 3.695000  1.915000 4.025000 2.635000 ;
      RECT 4.195000  0.255000 4.365000 0.615000 ;
      RECT 4.195000  0.615000 5.205000 0.785000 ;
      RECT 4.195000  1.935000 5.205000 2.105000 ;
      RECT 4.195000  2.105000 4.365000 2.465000 ;
      RECT 4.535000  0.085000 4.865000 0.445000 ;
      RECT 4.535000  2.275000 4.865000 2.635000 ;
      RECT 5.035000  0.255000 5.205000 0.615000 ;
      RECT 5.035000  2.105000 5.205000 2.465000 ;
      RECT 5.250000  0.955000 5.935000 1.125000 ;
      RECT 5.420000  0.765000 5.935000 0.955000 ;
      RECT 5.485000  2.125000 6.685000 2.465000 ;
      RECT 5.540000  0.255000 6.550000 0.505000 ;
      RECT 5.540000  0.505000 5.710000 0.595000 ;
      RECT 6.380000  0.505000 6.550000 0.655000 ;
      RECT 6.380000  0.655000 7.300000 0.825000 ;
      RECT 6.515000  1.935000 7.180000 2.105000 ;
      RECT 6.515000  2.105000 6.685000 2.125000 ;
      RECT 6.780000  0.085000 7.110000 0.445000 ;
      RECT 6.890000  2.275000 7.220000 2.635000 ;
      RECT 7.010000  1.470000 7.300000 1.640000 ;
      RECT 7.010000  1.640000 7.180000 1.935000 ;
      RECT 7.130000  0.825000 7.300000 1.075000 ;
      RECT 7.130000  1.075000 7.800000 1.245000 ;
      RECT 7.130000  1.245000 7.300000 1.470000 ;
      RECT 7.815000  1.795000 7.985000 2.635000 ;
      RECT 7.895000  0.085000 8.065000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  0.765000 2.155000 0.935000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.685000  0.765000 5.855000 0.935000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
    LAYER met1 ;
      RECT 1.925000 0.735000 2.215000 0.780000 ;
      RECT 1.925000 0.780000 5.915000 0.920000 ;
      RECT 1.925000 0.920000 2.215000 0.965000 ;
      RECT 5.625000 0.735000 5.915000 0.780000 ;
      RECT 5.625000 0.920000 5.915000 0.965000 ;
  END
END sky130_fd_sc_hd__fa_2
MACRO sky130_fd_sc_hd__fa_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fa_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.633000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.080000 0.995000 2.680000 1.275000 ;
        RECT 2.080000 1.275000 2.340000 1.325000 ;
      LAYER mcon ;
        RECT 2.450000 1.105000 2.620000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.610000 1.030000 4.000000 1.360000 ;
      LAYER mcon ;
        RECT 3.830000 1.105000 4.000000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.645000 0.955000 6.005000 1.275000 ;
      LAYER mcon ;
        RECT 5.690000 1.105000 5.860000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.030000 0.995000 7.885000 1.275000 ;
      LAYER mcon ;
        RECT 7.070000 1.105000 7.240000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.390000 1.075000 2.680000 1.120000 ;
        RECT 2.390000 1.120000 7.300000 1.260000 ;
        RECT 2.390000 1.260000 2.680000 1.305000 ;
        RECT 3.770000 1.075000 4.060000 1.120000 ;
        RECT 3.770000 1.260000 4.060000 1.305000 ;
        RECT 5.630000 1.075000 5.920000 1.120000 ;
        RECT 5.630000 1.260000 5.920000 1.305000 ;
        RECT 7.010000 1.075000 7.300000 1.120000 ;
        RECT 7.010000 1.260000 7.300000 1.305000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.633000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.480000 1.445000 3.080000 1.690000 ;
      LAYER mcon ;
        RECT 2.910000 1.445000 3.080000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.580000 1.435000 4.995000 1.745000 ;
      LAYER mcon ;
        RECT 4.770000 1.445000 4.940000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.075000 1.445000 7.760000 1.735000 ;
      LAYER mcon ;
        RECT 7.530000 1.445000 7.700000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.850000 1.415000 3.140000 1.460000 ;
        RECT 2.850000 1.460000 7.760000 1.600000 ;
        RECT 2.850000 1.600000 3.140000 1.645000 ;
        RECT 4.710000 1.415000 5.000000 1.460000 ;
        RECT 4.710000 1.600000 5.000000 1.645000 ;
        RECT 7.470000 1.415000 7.760000 1.460000 ;
        RECT 7.470000 1.600000 7.760000 1.645000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.477000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.050000 1.105000 3.420000 1.275000 ;
        RECT 3.250000 1.275000 3.420000 1.570000 ;
        RECT 3.250000 1.570000 4.340000 1.740000 ;
        RECT 4.170000 0.965000 5.390000 1.250000 ;
        RECT 4.170000 1.250000 4.340000 1.570000 ;
        RECT 5.220000 1.250000 5.390000 1.435000 ;
        RECT 5.220000 1.435000 5.580000 1.515000 ;
        RECT 5.220000 1.515000 6.845000 1.685000 ;
        RECT 6.595000 1.355000 6.845000 1.515000 ;
        RECT 6.595000 1.685000 6.845000 1.955000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.735000 1.525000 0.905000 ;
        RECT 0.085000 0.905000 0.435000 1.415000 ;
        RECT 0.085000 1.415000 1.570000 1.585000 ;
        RECT 0.515000 0.255000 0.845000 0.735000 ;
        RECT 0.515000 1.585000 0.845000 2.445000 ;
        RECT 1.355000 0.315000 1.685000 0.485000 ;
        RECT 1.355000 0.485000 1.525000 0.735000 ;
        RECT 1.400000 1.585000 1.570000 1.780000 ;
        RECT 1.400000 1.780000 1.645000 1.950000 ;
        RECT 1.435000 1.950000 1.645000 2.465000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.943000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.320000 0.255000  8.650000 0.485000 ;
        RECT 8.320000 1.795000  8.570000 1.965000 ;
        RECT 8.320000 1.965000  8.490000 2.465000 ;
        RECT 8.400000 0.485000  8.650000 0.735000 ;
        RECT 8.400000 0.735000 10.035000 0.905000 ;
        RECT 8.400000 1.415000 10.035000 1.585000 ;
        RECT 8.400000 1.585000  8.570000 1.795000 ;
        RECT 9.160000 0.270000  9.490000 0.735000 ;
        RECT 9.160000 1.585000  9.490000 2.425000 ;
        RECT 9.700000 0.905000 10.035000 1.415000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.175000  0.085000  0.345000 0.565000 ;
      RECT 0.175000  1.795000  0.345000 2.635000 ;
      RECT 0.605000  1.075000  1.910000 1.245000 ;
      RECT 1.015000  0.085000  1.185000 0.565000 ;
      RECT 1.015000  1.795000  1.185000 2.635000 ;
      RECT 1.740000  0.655000  3.090000 0.825000 ;
      RECT 1.740000  0.825000  1.910000 1.075000 ;
      RECT 1.740000  1.245000  1.910000 1.430000 ;
      RECT 1.740000  1.430000  1.945000 1.495000 ;
      RECT 1.740000  1.495000  2.310000 1.600000 ;
      RECT 1.775000  1.600000  2.310000 1.665000 ;
      RECT 1.815000  2.275000  2.145000 2.635000 ;
      RECT 1.855000  0.085000  2.185000 0.465000 ;
      RECT 2.140000  1.665000  2.310000 1.910000 ;
      RECT 2.140000  1.910000  3.170000 2.080000 ;
      RECT 2.370000  0.255000  3.090000 0.655000 ;
      RECT 2.735000  2.080000  3.170000 2.465000 ;
      RECT 2.850000  0.825000  3.090000 0.935000 ;
      RECT 3.340000  0.255000  3.510000 0.615000 ;
      RECT 3.340000  0.615000  4.350000 0.785000 ;
      RECT 3.340000  1.935000  4.415000 2.105000 ;
      RECT 3.340000  2.105000  3.510000 2.465000 ;
      RECT 3.680000  0.085000  4.010000 0.445000 ;
      RECT 3.680000  2.275000  4.010000 2.635000 ;
      RECT 4.180000  0.255000  4.350000 0.615000 ;
      RECT 4.180000  2.105000  4.415000 2.465000 ;
      RECT 4.620000  0.085000  4.950000 0.490000 ;
      RECT 4.620000  1.915000  4.950000 2.635000 ;
      RECT 5.120000  0.255000  5.290000 0.615000 ;
      RECT 5.120000  0.615000  6.130000 0.785000 ;
      RECT 5.120000  1.935000  6.130000 2.105000 ;
      RECT 5.120000  2.105000  5.290000 2.465000 ;
      RECT 5.460000  0.085000  5.790000 0.445000 ;
      RECT 5.460000  2.275000  5.790000 2.635000 ;
      RECT 5.960000  0.255000  6.130000 0.615000 ;
      RECT 5.960000  2.105000  6.130000 2.465000 ;
      RECT 6.175000  0.955000  6.860000 1.125000 ;
      RECT 6.345000  0.765000  6.860000 0.955000 ;
      RECT 6.410000  2.125000  7.610000 2.465000 ;
      RECT 6.465000  0.255000  7.475000 0.505000 ;
      RECT 6.465000  0.505000  6.635000 0.595000 ;
      RECT 7.305000  0.505000  7.475000 0.655000 ;
      RECT 7.305000  0.655000  8.225000 0.825000 ;
      RECT 7.440000  1.935000  8.105000 2.105000 ;
      RECT 7.440000  2.105000  7.610000 2.125000 ;
      RECT 7.705000  0.085000  8.035000 0.445000 ;
      RECT 7.815000  2.275000  8.145000 2.635000 ;
      RECT 7.935000  1.470000  8.225000 1.640000 ;
      RECT 7.935000  1.640000  8.105000 1.935000 ;
      RECT 8.055000  0.825000  8.225000 1.075000 ;
      RECT 8.055000  1.075000  9.445000 1.245000 ;
      RECT 8.055000  1.245000  8.225000 1.470000 ;
      RECT 8.740000  1.795000  8.910000 2.635000 ;
      RECT 8.820000  0.085000  8.990000 0.565000 ;
      RECT 9.660000  0.085000  9.830000 0.565000 ;
      RECT 9.660000  1.795000  9.830000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.910000  0.765000 3.080000 0.935000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.610000  0.765000 6.780000 0.935000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
    LAYER met1 ;
      RECT 2.850000 0.735000 3.140000 0.780000 ;
      RECT 2.850000 0.780000 6.840000 0.920000 ;
      RECT 2.850000 0.920000 3.140000 0.965000 ;
      RECT 6.550000 0.735000 6.840000 0.780000 ;
      RECT 6.550000 0.920000 6.840000 0.965000 ;
  END
END sky130_fd_sc_hd__fa_4
MACRO sky130_fd_sc_hd__fah_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fah_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.42000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 1.075000 1.440000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.691500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 1.075000 2.495000 1.275000 ;
        RECT 1.990000 1.275000 2.190000 1.410000 ;
        RECT 2.015000 1.410000 2.190000 1.725000 ;
      LAYER mcon ;
        RECT 1.990000 1.105000 2.160000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.675000 0.995000 5.925000 1.325000 ;
      LAYER mcon ;
        RECT 5.680000 1.105000 5.850000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.930000 1.075000 2.220000 1.120000 ;
        RECT 1.930000 1.120000 5.910000 1.260000 ;
        RECT 1.930000 1.260000 2.220000 1.305000 ;
        RECT 5.620000 1.075000 5.910000 1.120000 ;
        RECT 5.620000 1.260000 5.910000 1.305000 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.475000 1.075000  9.865000 1.325000 ;
        RECT 9.690000 0.735000 10.010000 0.935000 ;
        RECT 9.690000 0.935000  9.865000 1.075000 ;
    END
  END CI
  PIN COUT
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.870000 0.270000 11.310000 0.825000 ;
        RECT 10.870000 0.825000 11.040000 1.495000 ;
        RECT 10.870000 1.495000 11.390000 2.465000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.506000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.980000 0.255000 12.335000 0.825000 ;
        RECT 11.985000 1.785000 12.335000 2.465000 ;
        RECT 12.110000 0.825000 12.335000 1.785000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.420000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.610000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.420000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.420000 0.085000 ;
      RECT  0.000000  2.635000 12.420000 2.805000 ;
      RECT  0.085000  0.255000  0.425000 0.805000 ;
      RECT  0.085000  0.805000  0.255000 1.500000 ;
      RECT  0.085000  1.500000  0.445000 1.895000 ;
      RECT  0.085000  1.895000  2.805000 2.065000 ;
      RECT  0.085000  2.065000  0.395000 2.465000 ;
      RECT  0.425000  0.995000  0.780000 1.325000 ;
      RECT  0.565000  2.260000  0.930000 2.635000 ;
      RECT  0.595000  0.085000  0.765000 0.545000 ;
      RECT  0.595000  0.735000  1.320000 0.905000 ;
      RECT  0.595000  0.905000  0.780000 0.995000 ;
      RECT  0.610000  1.325000  0.780000 1.380000 ;
      RECT  0.610000  1.380000  0.815000 1.445000 ;
      RECT  0.610000  1.445000  1.315000 1.455000 ;
      RECT  0.615000  1.455000  1.315000 1.615000 ;
      RECT  0.985000  1.615000  1.315000 1.715000 ;
      RECT  0.990000  0.255000  1.320000 0.735000 ;
      RECT  1.490000  1.445000  1.820000 1.500000 ;
      RECT  1.490000  1.500000  1.840000 1.725000 ;
      RECT  1.500000  0.255000  1.840000 0.715000 ;
      RECT  1.500000  0.715000  2.520000 0.885000 ;
      RECT  1.500000  0.885000  1.820000 0.905000 ;
      RECT  1.615000  0.905000  1.820000 1.445000 ;
      RECT  2.010000  0.085000  2.180000 0.545000 ;
      RECT  2.065000  2.235000  2.395000 2.635000 ;
      RECT  2.350000  0.255000  4.840000 0.425000 ;
      RECT  2.350000  0.425000  2.520000 0.715000 ;
      RECT  2.360000  1.445000  2.860000 1.715000 ;
      RECT  2.635000  2.065000  2.805000 2.295000 ;
      RECT  2.635000  2.295000  4.950000 2.465000 ;
      RECT  2.690000  0.595000  2.860000 1.445000 ;
      RECT  3.030000  0.425000  4.840000 0.465000 ;
      RECT  3.030000  0.465000  3.200000 1.955000 ;
      RECT  3.030000  1.955000  4.320000 2.125000 ;
      RECT  3.370000  0.635000  3.900000 0.805000 ;
      RECT  3.370000  0.805000  3.540000 1.455000 ;
      RECT  3.370000  1.455000  3.815000 1.785000 ;
      RECT  3.985000  1.785000  4.320000 1.955000 ;
      RECT  4.070000  0.645000  4.400000 0.735000 ;
      RECT  4.070000  0.735000  4.560000 0.755000 ;
      RECT  4.070000  0.755000  5.170000 0.780000 ;
      RECT  4.070000  0.780000  5.155000 0.805000 ;
      RECT  4.070000  0.805000  5.145000 0.905000 ;
      RECT  4.070000  1.075000  4.400000 1.160000 ;
      RECT  4.070000  1.160000  4.535000 1.615000 ;
      RECT  4.480000  0.905000  5.145000 0.925000 ;
      RECT  4.650000  0.465000  4.840000 0.585000 ;
      RECT  4.705000  0.925000  4.875000 2.295000 ;
      RECT  4.925000  0.735000  5.180000 0.740000 ;
      RECT  4.925000  0.740000  5.170000 0.755000 ;
      RECT  4.950000  0.715000  5.180000 0.735000 ;
      RECT  4.980000  0.690000  5.180000 0.715000 ;
      RECT  5.000000  0.655000  5.180000 0.690000 ;
      RECT  5.010000  0.255000  6.100000 0.425000 ;
      RECT  5.010000  0.425000  5.180000 0.655000 ;
      RECT  5.125000  1.150000  5.505000 1.320000 ;
      RECT  5.125000  1.320000  5.295000 2.295000 ;
      RECT  5.125000  2.295000  7.560000 2.465000 ;
      RECT  5.320000  0.865000  5.520000 0.925000 ;
      RECT  5.320000  0.925000  5.505000 1.150000 ;
      RECT  5.335000  0.840000  5.520000 0.865000 ;
      RECT  5.350000  0.595000  5.520000 0.840000 ;
      RECT  5.475000  1.700000  5.875000 2.030000 ;
      RECT  5.750000  0.425000  6.100000 0.565000 ;
      RECT  6.105000  0.740000  6.435000 1.275000 ;
      RECT  6.105000  1.445000  6.460000 1.615000 ;
      RECT  6.270000  0.255000  9.735000 0.425000 ;
      RECT  6.270000  0.425000  6.600000 0.570000 ;
      RECT  6.290000  1.615000  6.460000 1.955000 ;
      RECT  6.290000  1.955000  7.220000 2.125000 ;
      RECT  6.610000  0.755000  6.940000 0.925000 ;
      RECT  6.610000  0.925000  6.880000 1.275000 ;
      RECT  6.710000  1.275000  6.880000 1.785000 ;
      RECT  6.770000  0.595000  6.940000 0.755000 ;
      RECT  7.050000  1.060000  7.280000 1.130000 ;
      RECT  7.050000  1.130000  7.245000 1.175000 ;
      RECT  7.050000  1.175000  7.220000 1.955000 ;
      RECT  7.065000  1.045000  7.280000 1.060000 ;
      RECT  7.090000  1.010000  7.280000 1.045000 ;
      RECT  7.110000  0.595000  7.445000 0.765000 ;
      RECT  7.110000  0.765000  7.280000 1.010000 ;
      RECT  7.390000  1.275000  7.620000 1.375000 ;
      RECT  7.390000  1.375000  7.595000 1.400000 ;
      RECT  7.390000  1.400000  7.575000 1.425000 ;
      RECT  7.390000  1.425000  7.560000 2.295000 ;
      RECT  7.450000  0.995000  7.620000 1.275000 ;
      RECT  7.705000  0.425000  7.960000 0.825000 ;
      RECT  7.730000  1.510000  7.960000 2.295000 ;
      RECT  7.730000  2.295000  9.655000 2.465000 ;
      RECT  7.790000  0.825000  7.960000 1.510000 ;
      RECT  8.145000  1.955000  9.250000 2.125000 ;
      RECT  8.155000  0.595000  8.405000 0.925000 ;
      RECT  8.225000  0.925000  8.405000 1.445000 ;
      RECT  8.225000  1.445000  8.910000 1.785000 ;
      RECT  8.575000  0.595000  8.745000 1.105000 ;
      RECT  8.575000  1.105000  9.250000 1.275000 ;
      RECT  8.920000  0.685000  9.300000 0.935000 ;
      RECT  9.080000  1.275000  9.250000 1.955000 ;
      RECT  9.400000  0.425000  9.735000 0.515000 ;
      RECT  9.420000  1.495000 10.350000 1.705000 ;
      RECT  9.420000  1.705000  9.655000 2.295000 ;
      RECT  9.840000  2.275000 10.175000 2.635000 ;
      RECT  9.905000  0.085000 10.075000 0.565000 ;
      RECT 10.180000  0.995000 10.350000 1.495000 ;
      RECT 10.245000  0.285000 10.690000 0.825000 ;
      RECT 10.345000  1.875000 10.690000 2.465000 ;
      RECT 10.520000  0.825000 10.690000 1.875000 ;
      RECT 11.210000  0.995000 11.460000 1.325000 ;
      RECT 11.480000  0.085000 11.810000 0.825000 ;
      RECT 11.560000  1.785000 11.815000 2.635000 ;
      RECT 11.630000  0.995000 11.940000 1.615000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.450000  1.445000  2.620000 1.615000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.370000  0.765000  3.540000 0.935000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.365000  1.445000  4.535000 1.615000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.570000  1.785000  5.740000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.150000  0.765000  6.320000 0.935000 ;
      RECT  6.150000  1.445000  6.320000 1.615000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.610000  1.105000  6.780000 1.275000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.460000  1.445000  8.630000 1.615000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  8.920000  0.765000  9.090000 0.935000 ;
      RECT  9.080000  1.785000  9.250000 1.955000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.520000  1.785000 10.690000 1.955000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.220000  1.105000 11.390000 1.275000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 11.680000  1.445000 11.850000 1.615000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
    LAYER met1 ;
      RECT  2.390000 1.415000  2.680000 1.460000 ;
      RECT  2.390000 1.460000  6.380000 1.600000 ;
      RECT  2.390000 1.600000  2.680000 1.645000 ;
      RECT  3.310000 0.735000  3.600000 0.780000 ;
      RECT  3.310000 0.780000  9.150000 0.920000 ;
      RECT  3.310000 0.920000  3.600000 0.965000 ;
      RECT  3.925000 1.755000  4.215000 1.800000 ;
      RECT  3.925000 1.800000  5.800000 1.940000 ;
      RECT  3.925000 1.940000  4.215000 1.985000 ;
      RECT  4.305000 1.415000  4.595000 1.460000 ;
      RECT  4.305000 1.600000  4.595000 1.645000 ;
      RECT  5.510000 1.755000  5.800000 1.800000 ;
      RECT  5.510000 1.940000  5.800000 1.985000 ;
      RECT  6.090000 0.735000  6.380000 0.780000 ;
      RECT  6.090000 0.920000  6.380000 0.965000 ;
      RECT  6.090000 1.415000  6.380000 1.460000 ;
      RECT  6.090000 1.600000  6.380000 1.645000 ;
      RECT  6.550000 1.075000  6.840000 1.120000 ;
      RECT  6.550000 1.120000 11.450000 1.260000 ;
      RECT  6.550000 1.260000  6.840000 1.305000 ;
      RECT  8.400000 1.415000  8.690000 1.460000 ;
      RECT  8.400000 1.460000 11.910000 1.600000 ;
      RECT  8.400000 1.600000  8.690000 1.645000 ;
      RECT  8.860000 0.735000  9.150000 0.780000 ;
      RECT  8.860000 0.920000  9.150000 0.965000 ;
      RECT  9.020000 1.755000  9.310000 1.800000 ;
      RECT  9.020000 1.800000 10.750000 1.940000 ;
      RECT  9.020000 1.940000  9.310000 1.985000 ;
      RECT 10.460000 1.755000 10.750000 1.800000 ;
      RECT 10.460000 1.940000 10.750000 1.985000 ;
      RECT 11.160000 1.075000 11.450000 1.120000 ;
      RECT 11.160000 1.260000 11.450000 1.305000 ;
      RECT 11.620000 1.415000 11.910000 1.460000 ;
      RECT 11.620000 1.600000 11.910000 1.645000 ;
  END
END sky130_fd_sc_hd__fah_1
MACRO sky130_fd_sc_hd__fahcin_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fahcin_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.42000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 1.075000 1.340000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.691500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.510000 0.665000 1.740000 1.325000 ;
      LAYER mcon ;
        RECT 1.525000 0.765000 1.695000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.240000 0.645000 4.490000 1.325000 ;
      LAYER mcon ;
        RECT 4.285000 0.765000 4.455000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465000 0.735000 1.755000 0.780000 ;
        RECT 1.465000 0.780000 4.515000 0.920000 ;
        RECT 1.465000 0.920000 1.755000 0.965000 ;
        RECT 4.225000 0.735000 4.515000 0.780000 ;
        RECT 4.225000 0.920000 4.515000 0.965000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.493500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.520000 1.075000 10.965000 1.275000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.402800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.600000 0.755000 6.925000 0.925000 ;
        RECT 6.600000 0.925000 6.870000 1.675000 ;
        RECT 6.700000 1.675000 6.870000 1.785000 ;
        RECT 6.755000 0.595000 6.925000 0.755000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.470250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.995000 0.255000 12.335000 0.825000 ;
        RECT 12.000000 1.785000 12.335000 2.465000 ;
        RECT 12.125000 0.825000 12.335000 1.785000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.420000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.610000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.420000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.420000 0.085000 ;
      RECT  0.000000  2.635000 12.420000 2.805000 ;
      RECT  0.085000  0.735000  0.430000 0.805000 ;
      RECT  0.085000  0.805000  0.255000 1.500000 ;
      RECT  0.085000  1.500000  0.440000 1.840000 ;
      RECT  0.085000  1.840000  1.110000 2.010000 ;
      RECT  0.085000  2.010000  0.430000 2.465000 ;
      RECT  0.100000  0.255000  0.430000 0.735000 ;
      RECT  0.425000  0.995000  0.780000 1.325000 ;
      RECT  0.600000  2.180000  0.770000 2.635000 ;
      RECT  0.610000  0.735000  1.325000 0.905000 ;
      RECT  0.610000  0.905000  0.780000 0.995000 ;
      RECT  0.610000  1.325000  0.780000 1.500000 ;
      RECT  0.610000  1.500000  1.450000 1.670000 ;
      RECT  0.630000  0.085000  0.800000 0.545000 ;
      RECT  0.940000  2.010000  1.110000 2.215000 ;
      RECT  0.940000  2.215000  1.970000 2.295000 ;
      RECT  0.940000  2.295000  3.515000 2.385000 ;
      RECT  0.995000  0.255000  3.390000 0.425000 ;
      RECT  0.995000  0.425000  2.100000 0.465000 ;
      RECT  0.995000  0.465000  1.325000 0.735000 ;
      RECT  1.280000  1.670000  1.450000 1.785000 ;
      RECT  1.280000  1.785000  2.050000 1.955000 ;
      RECT  1.280000  1.955000  1.450000 2.045000 ;
      RECT  1.715000  2.385000  3.515000 2.465000 ;
      RECT  1.985000  0.675000  2.390000 1.350000 ;
      RECT  2.220000  0.595000  2.390000 0.675000 ;
      RECT  2.220000  1.350000  2.390000 1.785000 ;
      RECT  2.515000  0.425000  3.390000 0.465000 ;
      RECT  2.565000  1.785000  2.895000 2.045000 ;
      RECT  2.620000  0.655000  3.025000 0.735000 ;
      RECT  2.620000  0.735000  3.135000 0.755000 ;
      RECT  2.620000  0.755000  3.730000 0.905000 ;
      RECT  2.640000  1.075000  2.970000 1.095000 ;
      RECT  2.640000  1.095000  3.120000 1.245000 ;
      RECT  2.800000  1.245000  3.120000 1.265000 ;
      RECT  2.950000  1.265000  3.120000 1.615000 ;
      RECT  3.055000  0.905000  3.730000 0.925000 ;
      RECT  3.215000  0.465000  3.390000 0.585000 ;
      RECT  3.245000  2.110000  3.460000 2.295000 ;
      RECT  3.290000  0.925000  3.460000 2.110000 ;
      RECT  3.560000  0.255000  4.570000 0.425000 ;
      RECT  3.560000  0.425000  3.730000 0.755000 ;
      RECT  3.710000  1.150000  4.070000 1.320000 ;
      RECT  3.710000  1.320000  3.880000 2.290000 ;
      RECT  3.710000  2.290000  5.065000 2.460000 ;
      RECT  3.900000  0.595000  4.070000 1.150000 ;
      RECT  4.080000  1.695000  4.445000 2.120000 ;
      RECT  4.240000  0.425000  4.570000 0.475000 ;
      RECT  4.690000  1.385000  5.170000 1.725000 ;
      RECT  4.815000  1.895000  5.995000 2.065000 ;
      RECT  4.815000  2.065000  5.065000 2.290000 ;
      RECT  4.830000  0.510000  5.000000 0.995000 ;
      RECT  4.830000  0.995000  5.630000 1.325000 ;
      RECT  4.830000  1.325000  5.170000 1.385000 ;
      RECT  5.180000  0.085000  5.510000 0.805000 ;
      RECT  5.260000  2.235000  5.590000 2.635000 ;
      RECT  5.635000  1.555000  6.370000 1.725000 ;
      RECT  5.680000  0.380000  5.970000 0.815000 ;
      RECT  5.800000  0.815000  5.970000 1.555000 ;
      RECT  5.825000  2.065000  5.995000 2.295000 ;
      RECT  5.825000  2.295000  7.950000 2.465000 ;
      RECT  6.140000  0.740000  6.425000 1.325000 ;
      RECT  6.200000  1.725000  6.370000 1.895000 ;
      RECT  6.200000  1.895000  6.530000 1.955000 ;
      RECT  6.200000  1.955000  7.210000 2.125000 ;
      RECT  6.255000  0.255000  7.695000 0.425000 ;
      RECT  6.255000  0.425000  6.585000 0.570000 ;
      RECT  7.040000  1.060000  7.270000 1.230000 ;
      RECT  7.040000  1.230000  7.210000 1.955000 ;
      RECT  7.100000  0.595000  7.350000 0.925000 ;
      RECT  7.100000  0.925000  7.270000 1.060000 ;
      RECT  7.380000  1.360000  7.610000 1.530000 ;
      RECT  7.380000  1.530000  7.550000 2.125000 ;
      RECT  7.440000  1.105000  7.695000 1.290000 ;
      RECT  7.440000  1.290000  7.610000 1.360000 ;
      RECT  7.520000  0.425000  7.695000 1.105000 ;
      RECT  7.780000  1.550000  8.035000 1.720000 ;
      RECT  7.780000  1.720000  7.950000 2.295000 ;
      RECT  7.865000  0.255000  9.980000 0.425000 ;
      RECT  7.865000  0.425000  8.035000 0.740000 ;
      RECT  7.865000  0.995000  8.035000 1.550000 ;
      RECT  8.220000  1.955000  8.390000 2.295000 ;
      RECT  8.220000  2.295000  9.410000 2.465000 ;
      RECT  8.305000  0.595000  8.555000 0.925000 ;
      RECT  8.375000  0.925000  8.555000 1.445000 ;
      RECT  8.375000  1.445000  8.670000 1.530000 ;
      RECT  8.375000  1.530000  8.890000 1.785000 ;
      RECT  8.560000  1.785000  8.890000 2.125000 ;
      RECT  8.725000  0.595000  9.410000 0.765000 ;
      RECT  8.835000  0.995000  9.070000 1.325000 ;
      RECT  9.240000  0.765000  9.410000 1.875000 ;
      RECT  9.240000  1.875000 10.885000 2.025000 ;
      RECT  9.240000  2.025000 10.145000 2.030000 ;
      RECT  9.240000  2.030000 10.130000 2.035000 ;
      RECT  9.240000  2.035000 10.120000 2.040000 ;
      RECT  9.240000  2.040000 10.105000 2.045000 ;
      RECT  9.240000  2.045000  9.410000 2.295000 ;
      RECT  9.640000  0.425000  9.980000 0.825000 ;
      RECT  9.640000  0.825000  9.810000 1.535000 ;
      RECT  9.640000  1.535000 10.010000 1.705000 ;
      RECT  9.980000  0.995000 10.350000 1.325000 ;
      RECT 10.055000  1.870000 10.885000 1.875000 ;
      RECT 10.070000  1.865000 10.885000 1.870000 ;
      RECT 10.085000  1.860000 10.885000 1.865000 ;
      RECT 10.100000  1.855000 10.885000 1.860000 ;
      RECT 10.180000  0.085000 10.350000 0.565000 ;
      RECT 10.180000  0.735000 10.910000 0.905000 ;
      RECT 10.180000  0.905000 10.350000 0.995000 ;
      RECT 10.180000  1.325000 10.350000 1.445000 ;
      RECT 10.180000  1.445000 10.885000 1.855000 ;
      RECT 10.190000  2.195000 10.360000 2.635000 ;
      RECT 10.530000  0.285000 10.910000 0.735000 ;
      RECT 10.535000  2.025000 10.885000 2.465000 ;
      RECT 11.075000  1.455000 11.405000 2.465000 ;
      RECT 11.155000  0.270000 11.325000 0.680000 ;
      RECT 11.155000  0.680000 11.405000 1.455000 ;
      RECT 11.495000  0.085000 11.825000 0.510000 ;
      RECT 11.575000  1.785000 11.830000 2.635000 ;
      RECT 11.645000  0.995000 11.955000 1.615000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.880000  1.785000  2.050000 1.955000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  1.105000  2.155000 1.275000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.570000  1.785000  2.740000 1.955000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  2.950000  1.445000  3.120000 1.615000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.140000  1.785000  4.310000 1.955000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.760000  1.445000  4.930000 1.615000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.140000  1.105000  6.310000 1.275000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.520000  0.765000  7.690000 0.935000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.440000  1.445000  8.610000 1.615000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  8.900000  1.105000  9.070000 1.275000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.220000  0.765000 11.390000 0.935000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 11.680000  1.445000 11.850000 1.615000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
    LAYER met1 ;
      RECT  1.820000 1.755000  2.110000 1.800000 ;
      RECT  1.820000 1.800000  4.370000 1.940000 ;
      RECT  1.820000 1.940000  2.110000 1.985000 ;
      RECT  1.925000 1.075000  2.215000 1.120000 ;
      RECT  1.925000 1.120000  9.130000 1.260000 ;
      RECT  1.925000 1.260000  2.215000 1.305000 ;
      RECT  2.510000 1.755000  2.800000 1.800000 ;
      RECT  2.510000 1.940000  2.800000 1.985000 ;
      RECT  2.890000 1.415000  3.180000 1.460000 ;
      RECT  2.890000 1.460000  4.990000 1.600000 ;
      RECT  2.890000 1.600000  3.180000 1.645000 ;
      RECT  4.080000 1.755000  4.370000 1.800000 ;
      RECT  4.080000 1.940000  4.370000 1.985000 ;
      RECT  4.700000 1.415000  4.990000 1.460000 ;
      RECT  4.700000 1.600000  4.990000 1.645000 ;
      RECT  6.080000 1.075000  6.370000 1.120000 ;
      RECT  6.080000 1.260000  6.370000 1.305000 ;
      RECT  7.460000 0.735000  7.750000 0.780000 ;
      RECT  7.460000 0.780000 11.450000 0.920000 ;
      RECT  7.460000 0.920000  7.750000 0.965000 ;
      RECT  8.380000 1.415000  8.670000 1.460000 ;
      RECT  8.380000 1.460000 11.910000 1.600000 ;
      RECT  8.380000 1.600000  8.670000 1.645000 ;
      RECT  8.840000 1.075000  9.130000 1.120000 ;
      RECT  8.840000 1.260000  9.130000 1.305000 ;
      RECT 11.160000 0.735000 11.450000 0.780000 ;
      RECT 11.160000 0.920000 11.450000 0.965000 ;
      RECT 11.620000 1.415000 11.910000 1.460000 ;
      RECT 11.620000 1.600000 11.910000 1.645000 ;
  END
END sky130_fd_sc_hd__fahcin_1
MACRO sky130_fd_sc_hd__fahcon_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fahcon_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.42000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 1.075000 1.340000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.937500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.510000 0.710000 1.780000 1.325000 ;
      LAYER mcon ;
        RECT 1.525000 0.765000 1.695000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.265000 0.645000 4.515000 1.325000 ;
      LAYER mcon ;
        RECT 4.310000 0.765000 4.480000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465000 0.735000 1.755000 0.780000 ;
        RECT 1.465000 0.780000 4.540000 0.920000 ;
        RECT 1.465000 0.920000 1.755000 0.965000 ;
        RECT 4.250000 0.735000 4.540000 0.780000 ;
        RECT 4.250000 0.920000 4.540000 0.965000 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.493500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.530000 1.075000 10.975000 1.275000 ;
    END
  END CI
  PIN COUT_N
    ANTENNADIFFAREA  0.402800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.610000 0.755000 6.935000 0.925000 ;
        RECT 6.610000 0.925000 6.880000 1.675000 ;
        RECT 6.710000 1.675000 6.880000 1.785000 ;
        RECT 6.765000 0.595000 6.935000 0.755000 ;
    END
  END COUT_N
  PIN SUM
    ANTENNADIFFAREA  0.463750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.995000 0.255000 12.335000 0.825000 ;
        RECT 12.010000 1.785000 12.335000 2.465000 ;
        RECT 12.135000 0.825000 12.335000 1.785000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.420000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.610000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.420000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.420000 0.085000 ;
      RECT  0.000000  2.635000 12.420000 2.805000 ;
      RECT  0.085000  0.735000  0.430000 0.805000 ;
      RECT  0.085000  0.805000  0.255000 1.500000 ;
      RECT  0.085000  1.500000  0.440000 1.840000 ;
      RECT  0.085000  1.840000  1.110000 2.010000 ;
      RECT  0.085000  2.010000  0.430000 2.465000 ;
      RECT  0.100000  0.255000  0.430000 0.735000 ;
      RECT  0.425000  0.995000  0.780000 1.325000 ;
      RECT  0.600000  2.180000  0.770000 2.635000 ;
      RECT  0.610000  0.735000  1.325000 0.905000 ;
      RECT  0.610000  0.905000  0.780000 0.995000 ;
      RECT  0.610000  1.325000  0.780000 1.500000 ;
      RECT  0.610000  1.500000  1.450000 1.670000 ;
      RECT  0.630000  0.085000  0.800000 0.545000 ;
      RECT  0.940000  2.010000  1.110000 2.215000 ;
      RECT  0.940000  2.215000  2.545000 2.295000 ;
      RECT  0.940000  2.295000  3.540000 2.385000 ;
      RECT  0.995000  0.255000  3.410000 0.465000 ;
      RECT  0.995000  0.465000  1.325000 0.735000 ;
      RECT  1.280000  1.670000  1.450000 1.875000 ;
      RECT  1.280000  1.875000  2.920000 2.045000 ;
      RECT  1.965000  0.635000  2.470000 1.705000 ;
      RECT  2.375000  2.385000  3.540000 2.465000 ;
      RECT  2.640000  0.655000  3.025000 0.735000 ;
      RECT  2.640000  0.735000  3.160000 0.755000 ;
      RECT  2.640000  0.755000  3.750000 0.905000 ;
      RECT  2.640000  1.075000  2.975000 1.160000 ;
      RECT  2.640000  1.160000  3.100000 1.615000 ;
      RECT  3.055000  0.905000  3.750000 0.925000 ;
      RECT  3.240000  0.465000  3.410000 0.585000 ;
      RECT  3.270000  0.925000  3.440000 2.295000 ;
      RECT  3.580000  0.255000  4.595000 0.425000 ;
      RECT  3.580000  0.425000  3.750000 0.755000 ;
      RECT  3.725000  1.150000  4.095000 1.320000 ;
      RECT  3.725000  1.320000  3.895000 2.295000 ;
      RECT  3.725000  2.295000  5.100000 2.465000 ;
      RECT  3.925000  0.595000  4.095000 1.150000 ;
      RECT  4.210000  1.755000  4.380000 2.095000 ;
      RECT  4.265000  0.425000  4.595000 0.475000 ;
      RECT  4.700000  1.385000  5.180000 1.725000 ;
      RECT  4.840000  0.510000  5.030000 0.995000 ;
      RECT  4.840000  0.995000  5.180000 1.385000 ;
      RECT  4.875000  1.895000  6.005000 2.065000 ;
      RECT  4.875000  2.065000  5.100000 2.295000 ;
      RECT  5.200000  0.085000  5.530000 0.805000 ;
      RECT  5.270000  2.235000  5.600000 2.635000 ;
      RECT  5.645000  1.555000  6.380000 1.725000 ;
      RECT  5.700000  0.380000  5.980000 0.815000 ;
      RECT  5.810000  0.815000  5.980000 1.555000 ;
      RECT  5.835000  2.065000  6.005000 2.295000 ;
      RECT  5.835000  2.295000  7.960000 2.465000 ;
      RECT  6.150000  0.740000  6.435000 1.325000 ;
      RECT  6.210000  1.725000  6.380000 1.895000 ;
      RECT  6.210000  1.895000  6.540000 1.955000 ;
      RECT  6.210000  1.955000  7.220000 2.125000 ;
      RECT  6.265000  0.255000  7.700000 0.425000 ;
      RECT  6.265000  0.425000  6.595000 0.570000 ;
      RECT  7.050000  1.060000  7.280000 1.230000 ;
      RECT  7.050000  1.230000  7.220000 1.955000 ;
      RECT  7.110000  0.595000  7.360000 0.925000 ;
      RECT  7.110000  0.925000  7.280000 1.060000 ;
      RECT  7.390000  1.360000  7.620000 1.530000 ;
      RECT  7.390000  1.530000  7.560000 2.125000 ;
      RECT  7.450000  1.105000  7.700000 1.290000 ;
      RECT  7.450000  1.290000  7.620000 1.360000 ;
      RECT  7.530000  0.425000  7.700000 1.105000 ;
      RECT  7.790000  1.550000  8.045000 1.720000 ;
      RECT  7.790000  1.720000  7.960000 2.295000 ;
      RECT  7.875000  0.995000  8.045000 1.550000 ;
      RECT  7.935000  0.255000  9.450000 0.425000 ;
      RECT  7.935000  0.425000  8.270000 0.825000 ;
      RECT  8.230000  1.785000  8.400000 2.295000 ;
      RECT  8.230000  2.295000  9.950000 2.465000 ;
      RECT  8.440000  0.595000  8.900000 0.765000 ;
      RECT  8.440000  0.765000  8.610000 1.445000 ;
      RECT  8.440000  1.445000  8.740000 1.530000 ;
      RECT  8.440000  1.530000  8.900000 1.615000 ;
      RECT  8.570000  1.615000  8.900000 2.125000 ;
      RECT  8.780000  0.995000  9.110000 1.275000 ;
      RECT  9.070000  1.530000  9.450000 2.045000 ;
      RECT  9.070000  2.045000  9.420000 2.125000 ;
      RECT  9.280000  0.425000  9.450000 1.530000 ;
      RECT  9.620000  2.215000  9.950000 2.295000 ;
      RECT  9.650000  0.255000 10.020000 0.825000 ;
      RECT  9.650000  0.825000  9.820000 1.535000 ;
      RECT  9.650000  1.535000  9.950000 2.215000 ;
      RECT  9.990000  0.995000 10.360000 1.325000 ;
      RECT 10.120000  2.275000 10.455000 2.635000 ;
      RECT 10.190000  0.735000 10.920000 0.905000 ;
      RECT 10.190000  0.905000 10.360000 0.995000 ;
      RECT 10.190000  1.325000 10.360000 1.455000 ;
      RECT 10.190000  1.455000 10.835000 2.045000 ;
      RECT 10.200000  0.085000 10.370000 0.565000 ;
      RECT 10.540000  0.285000 10.920000 0.735000 ;
      RECT 10.625000  2.045000 10.835000 2.465000 ;
      RECT 11.085000  1.455000 11.415000 2.465000 ;
      RECT 11.165000  0.270000 11.335000 0.680000 ;
      RECT 11.165000  0.680000 11.415000 1.455000 ;
      RECT 11.535000  0.085000 11.825000 0.555000 ;
      RECT 11.585000  1.785000 11.840000 2.635000 ;
      RECT 11.655000  0.995000 11.965000 1.615000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.280000  1.785000  1.450000 1.955000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  1.105000  2.155000 1.275000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  2.930000  1.445000  3.100000 1.615000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.210000  1.785000  4.380000 1.955000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.770000  1.445000  4.940000 1.615000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.150000  1.105000  6.320000 1.275000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.530000  0.765000  7.700000 0.935000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.450000  1.445000  8.620000 1.615000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  8.910000  1.105000  9.080000 1.275000 ;
      RECT  9.280000  1.785000  9.450000 1.955000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.190000  1.785000 10.360000 1.955000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.230000  0.765000 11.400000 0.935000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 11.690000  1.445000 11.860000 1.615000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
    LAYER met1 ;
      RECT  1.195000 1.755000  1.510000 1.800000 ;
      RECT  1.195000 1.800000  4.440000 1.940000 ;
      RECT  1.195000 1.940000  1.510000 1.985000 ;
      RECT  1.925000 1.075000  2.215000 1.120000 ;
      RECT  1.925000 1.120000  9.140000 1.260000 ;
      RECT  1.925000 1.260000  2.215000 1.305000 ;
      RECT  2.845000 1.415000  3.160000 1.460000 ;
      RECT  2.845000 1.460000  5.000000 1.600000 ;
      RECT  2.845000 1.600000  3.160000 1.645000 ;
      RECT  4.150000 1.755000  4.440000 1.800000 ;
      RECT  4.150000 1.940000  4.440000 1.985000 ;
      RECT  4.710000 1.415000  5.000000 1.460000 ;
      RECT  4.710000 1.600000  5.000000 1.645000 ;
      RECT  6.090000 1.075000  6.380000 1.120000 ;
      RECT  6.090000 1.260000  6.380000 1.305000 ;
      RECT  7.470000 0.735000  7.760000 0.780000 ;
      RECT  7.470000 0.780000 11.460000 0.920000 ;
      RECT  7.470000 0.920000  7.760000 0.965000 ;
      RECT  8.390000 1.415000  8.680000 1.460000 ;
      RECT  8.390000 1.460000 11.920000 1.600000 ;
      RECT  8.390000 1.600000  8.680000 1.645000 ;
      RECT  8.850000 1.075000  9.140000 1.120000 ;
      RECT  8.850000 1.260000  9.140000 1.305000 ;
      RECT  9.195000 1.755000  9.510000 1.800000 ;
      RECT  9.195000 1.800000 10.420000 1.940000 ;
      RECT  9.195000 1.940000  9.510000 1.985000 ;
      RECT 10.130000 1.755000 10.420000 1.800000 ;
      RECT 10.130000 1.940000 10.420000 1.985000 ;
      RECT 11.170000 0.735000 11.460000 0.780000 ;
      RECT 11.170000 0.920000 11.460000 0.965000 ;
      RECT 11.630000 1.415000 11.920000 1.460000 ;
      RECT 11.630000 1.600000 11.920000 1.645000 ;
  END
END sky130_fd_sc_hd__fahcon_1
MACRO sky130_fd_sc_hd__fill_1
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.055000 0.260000 0.055000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
END sky130_fd_sc_hd__fill_1
MACRO sky130_fd_sc_hd__fill_2
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.920000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.920000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155000 -0.050000 0.315000 0.060000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.110000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.920000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.920000 0.085000 ;
      RECT 0.000000  2.635000 0.920000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
  END
END sky130_fd_sc_hd__fill_2
MACRO sky130_fd_sc_hd__fill_4
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.175000 -0.060000 0.285000 0.060000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__fill_4
MACRO sky130_fd_sc_hd__fill_8
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.130000 -0.120000 0.350000 0.050000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__fill_8
MACRO sky130_fd_sc_hd__ha_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ha_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335000 1.315000 3.585000 1.485000 ;
        RECT 3.360000 1.055000 3.585000 1.315000 ;
        RECT 3.360000 1.485000 3.585000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.850000 1.345000 2.155000 1.655000 ;
        RECT 1.850000 1.655000 3.165000 1.825000 ;
        RECT 1.850000 1.825000 2.155000 2.375000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175000 0.315000 4.515000 0.825000 ;
        RECT 4.175000 1.565000 4.515000 2.415000 ;
        RECT 4.330000 0.825000 4.515000 1.565000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.315000 0.425000 0.825000 ;
        RECT 0.090000 0.825000 0.320000 1.565000 ;
        RECT 0.090000 1.565000 0.425000 2.415000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.490000  1.075000 1.130000 1.245000 ;
      RECT 0.595000  0.085000 0.790000 0.885000 ;
      RECT 0.595000  1.515000 0.790000 2.275000 ;
      RECT 0.595000  2.275000 1.260000 2.635000 ;
      RECT 0.960000  0.345000 1.285000 0.675000 ;
      RECT 0.960000  0.675000 1.130000 1.075000 ;
      RECT 0.960000  1.245000 1.130000 1.935000 ;
      RECT 0.960000  1.935000 1.680000 2.105000 ;
      RECT 1.300000  0.975000 3.170000 1.145000 ;
      RECT 1.300000  1.145000 1.470000 1.325000 ;
      RECT 1.510000  2.105000 1.680000 2.355000 ;
      RECT 1.535000  0.345000 1.705000 0.635000 ;
      RECT 1.535000  0.635000 2.545000 0.805000 ;
      RECT 1.875000  0.085000 2.205000 0.465000 ;
      RECT 2.375000  0.345000 2.545000 0.635000 ;
      RECT 2.450000  2.275000 3.120000 2.635000 ;
      RECT 3.000000  0.345000 3.170000 0.715000 ;
      RECT 3.000000  0.715000 4.005000 0.885000 ;
      RECT 3.000000  0.885000 3.170000 0.975000 ;
      RECT 3.350000  1.785000 4.005000 1.955000 ;
      RECT 3.350000  1.955000 3.520000 2.355000 ;
      RECT 3.755000  0.085000 4.005000 0.545000 ;
      RECT 3.755000  2.125000 4.005000 2.635000 ;
      RECT 3.835000  0.885000 4.005000 0.995000 ;
      RECT 3.835000  0.995000 4.160000 1.325000 ;
      RECT 3.835000  1.325000 4.005000 1.785000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__ha_1
MACRO sky130_fd_sc_hd__ha_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ha_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 1.055000 4.045000 1.225000 ;
        RECT 3.820000 1.225000 4.045000 1.675000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.310000 1.005000 2.615000 1.395000 ;
        RECT 2.310000 1.395000 3.595000 1.675000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.635000 0.315000 4.965000 0.825000 ;
        RECT 4.715000 1.545000 4.965000 2.415000 ;
        RECT 4.790000 0.825000 4.965000 1.545000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 0.315000 0.885000 0.825000 ;
        RECT 0.555000 0.825000 0.780000 1.565000 ;
        RECT 0.555000 1.565000 0.885000 2.415000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.135000  0.085000 0.375000 0.885000 ;
      RECT 0.135000  1.495000 0.375000 2.635000 ;
      RECT 0.950000  1.075000 1.590000 1.245000 ;
      RECT 1.055000  0.085000 1.250000 0.885000 ;
      RECT 1.055000  1.515000 1.250000 2.635000 ;
      RECT 1.420000  0.345000 1.745000 0.675000 ;
      RECT 1.420000  0.675000 1.590000 1.075000 ;
      RECT 1.420000  1.245000 1.590000 2.205000 ;
      RECT 1.420000  2.205000 2.220000 2.375000 ;
      RECT 1.760000  0.995000 1.930000 1.855000 ;
      RECT 1.760000  1.855000 4.465000 2.025000 ;
      RECT 1.995000  0.345000 2.165000 0.635000 ;
      RECT 1.995000  0.635000 3.005000 0.805000 ;
      RECT 2.335000  0.085000 2.665000 0.465000 ;
      RECT 2.835000  0.345000 3.005000 0.635000 ;
      RECT 2.850000  2.205000 3.640000 2.635000 ;
      RECT 3.460000  0.345000 3.630000 0.715000 ;
      RECT 3.460000  0.715000 4.465000 0.885000 ;
      RECT 3.810000  2.025000 3.980000 2.355000 ;
      RECT 4.215000  0.085000 4.465000 0.545000 ;
      RECT 4.215000  2.205000 4.545000 2.635000 ;
      RECT 4.295000  0.885000 4.465000 0.995000 ;
      RECT 4.295000  0.995000 4.620000 1.325000 ;
      RECT 4.295000  1.325000 4.465000 1.855000 ;
      RECT 5.145000  0.085000 5.385000 0.885000 ;
      RECT 5.145000  1.495000 5.385000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__ha_2
MACRO sky130_fd_sc_hd__ha_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ha_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.320000 1.075000 4.380000 1.245000 ;
        RECT 4.210000 1.245000 4.380000 1.505000 ;
        RECT 4.210000 1.505000 6.810000 1.675000 ;
        RECT 5.625000 0.995000 5.795000 1.505000 ;
        RECT 6.580000 0.995000 7.055000 1.325000 ;
        RECT 6.580000 1.325000 6.810000 1.505000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.550000 0.995000 5.455000 1.165000 ;
        RECT 4.550000 1.165000 4.720000 1.325000 ;
        RECT 5.285000 0.730000 6.315000 0.825000 ;
        RECT 5.285000 0.825000 5.535000 0.845000 ;
        RECT 5.285000 0.845000 5.495000 0.875000 ;
        RECT 5.285000 0.875000 5.455000 0.995000 ;
        RECT 5.295000 0.720000 6.315000 0.730000 ;
        RECT 5.310000 0.710000 6.315000 0.720000 ;
        RECT 5.320000 0.695000 6.315000 0.710000 ;
        RECT 5.335000 0.675000 6.315000 0.695000 ;
        RECT 5.345000 0.655000 6.315000 0.675000 ;
        RECT 6.085000 0.825000 6.315000 1.325000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.595000 0.315000 7.845000 0.735000 ;
        RECT 7.595000 0.735000 8.685000 0.905000 ;
        RECT 7.595000 1.415000 8.685000 1.585000 ;
        RECT 7.595000 1.585000 7.765000 2.415000 ;
        RECT 8.405000 0.315000 8.685000 0.735000 ;
        RECT 8.405000 0.905000 8.685000 1.415000 ;
        RECT 8.405000 1.585000 8.685000 2.415000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.315000 0.845000 1.065000 ;
        RECT 0.515000 1.065000 1.550000 1.335000 ;
        RECT 0.515000 1.335000 0.845000 2.415000 ;
        RECT 1.355000 0.315000 1.685000 0.825000 ;
        RECT 1.355000 0.825000 1.550000 1.065000 ;
        RECT 1.355000 1.335000 1.550000 1.565000 ;
        RECT 1.355000 1.565000 1.685000 2.415000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.135000  0.085000 0.345000 0.885000 ;
      RECT 0.135000  1.495000 0.345000 2.635000 ;
      RECT 1.015000  0.085000 1.185000 0.885000 ;
      RECT 1.015000  1.515000 1.185000 2.635000 ;
      RECT 1.720000  1.075000 2.750000 1.245000 ;
      RECT 1.855000  0.085000 2.095000 0.885000 ;
      RECT 1.855000  1.495000 2.365000 2.635000 ;
      RECT 2.270000  0.305000 3.385000 0.475000 ;
      RECT 2.580000  0.645000 3.045000 0.815000 ;
      RECT 2.580000  0.815000 2.750000 1.075000 ;
      RECT 2.580000  1.245000 2.750000 1.765000 ;
      RECT 2.580000  1.765000 3.700000 1.935000 ;
      RECT 2.770000  1.935000 2.940000 2.355000 ;
      RECT 2.920000  0.995000 3.090000 1.425000 ;
      RECT 2.920000  1.425000 4.040000 1.595000 ;
      RECT 3.190000  2.105000 3.360000 2.635000 ;
      RECT 3.215000  0.475000 3.385000 0.645000 ;
      RECT 3.215000  0.645000 5.115000 0.815000 ;
      RECT 3.530000  1.935000 3.700000 2.205000 ;
      RECT 3.530000  2.205000 4.330000 2.375000 ;
      RECT 3.555000  0.085000 3.910000 0.465000 ;
      RECT 3.870000  1.595000 4.040000 1.855000 ;
      RECT 3.870000  1.855000 7.395000 2.025000 ;
      RECT 4.080000  0.345000 4.250000 0.645000 ;
      RECT 4.420000  0.085000 4.750000 0.465000 ;
      RECT 4.920000  0.255000 5.190000 0.585000 ;
      RECT 4.920000  0.585000 5.115000 0.645000 ;
      RECT 5.240000  2.205000 5.570000 2.635000 ;
      RECT 5.385000  0.085000 5.715000 0.465000 ;
      RECT 5.835000  2.025000 6.005000 2.355000 ;
      RECT 6.175000  0.295000 6.875000 0.465000 ;
      RECT 6.175000  2.205000 6.505000 2.635000 ;
      RECT 6.675000  2.025000 6.845000 2.355000 ;
      RECT 6.705000  0.465000 6.875000 0.645000 ;
      RECT 6.705000  0.645000 7.395000 0.815000 ;
      RECT 7.055000  0.085000 7.385000 0.465000 ;
      RECT 7.055000  2.205000 7.385000 2.635000 ;
      RECT 7.225000  0.815000 7.395000 1.075000 ;
      RECT 7.225000  1.075000 8.225000 1.245000 ;
      RECT 7.225000  1.245000 7.395000 1.855000 ;
      RECT 7.935000  1.755000 8.225000 2.635000 ;
      RECT 8.015000  0.085000 8.225000 0.565000 ;
      RECT 8.855000  0.085000 9.065000 0.885000 ;
      RECT 8.855000  1.495000 9.065000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
  END
END sky130_fd_sc_hd__ha_4
MACRO sky130_fd_sc_hd__inv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.320000 1.075000 0.650000 1.315000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.720000 0.255000 1.050000 0.885000 ;
        RECT 0.720000 1.485000 1.050000 2.465000 ;
        RECT 0.820000 0.885000 1.050000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.320000  0.085000 0.550000 0.905000 ;
      RECT 0.340000  1.495000 0.550000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__inv_1
MACRO sky130_fd_sc_hd__inv_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 0.435000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 0.255000 0.855000 0.885000 ;
        RECT 0.525000 1.485000 0.855000 2.465000 ;
        RECT 0.605000 0.885000 0.855000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.125000  0.085000 0.355000 0.905000 ;
      RECT 0.125000  1.495000 0.355000 2.635000 ;
      RECT 1.025000  0.085000 1.235000 0.905000 ;
      RECT 1.025000  1.495000 1.235000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__inv_2
MACRO sky130_fd_sc_hd__inv_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 1.735000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 0.255000 0.895000 0.725000 ;
        RECT 0.565000 0.725000 2.170000 0.905000 ;
        RECT 0.565000 1.495000 2.170000 1.665000 ;
        RECT 0.565000 1.665000 0.895000 2.465000 ;
        RECT 1.405000 0.255000 1.735000 0.725000 ;
        RECT 1.405000 1.665000 2.170000 1.685000 ;
        RECT 1.405000 1.685000 1.735000 2.465000 ;
        RECT 1.905000 0.905000 2.170000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.130000  0.085000 0.395000 0.545000 ;
      RECT 0.130000  1.495000 0.395000 2.635000 ;
      RECT 1.065000  0.085000 1.235000 0.545000 ;
      RECT 1.065000  1.835000 1.235000 2.635000 ;
      RECT 1.905000  0.085000 2.155000 0.550000 ;
      RECT 1.905000  2.175000 2.115000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__inv_4
MACRO sky130_fd_sc_hd__inv_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_6 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.485000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 2.615000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.336500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.685000 1.495000 3.135000 1.665000 ;
        RECT 0.685000 1.665000 1.015000 2.465000 ;
        RECT 0.765000 0.255000 0.935000 0.725000 ;
        RECT 0.765000 0.725000 3.135000 0.905000 ;
        RECT 1.525000 1.665000 1.855000 2.465000 ;
        RECT 1.605000 0.255000 1.775000 0.725000 ;
        RECT 2.365000 1.665000 3.135000 1.685000 ;
        RECT 2.365000 1.685000 2.695000 2.465000 ;
        RECT 2.445000 0.255000 2.615000 0.725000 ;
        RECT 2.785000 0.905000 3.135000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.130000  0.085000 0.395000 0.545000 ;
      RECT 0.130000  1.495000 0.425000 2.635000 ;
      RECT 1.185000  0.085000 1.355000 0.545000 ;
      RECT 1.185000  1.835000 1.355000 2.635000 ;
      RECT 2.025000  0.085000 2.195000 0.545000 ;
      RECT 2.025000  1.835000 2.195000 2.635000 ;
      RECT 2.785000  0.085000 3.035000 0.550000 ;
      RECT 2.865000  2.175000 3.035000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__inv_6
MACRO sky130_fd_sc_hd__inv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.680000 1.075000 3.535000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 4.055000 0.905000 ;
        RECT 0.085000 0.905000 0.430000 1.495000 ;
        RECT 0.085000 1.495000 4.055000 1.665000 ;
        RECT 0.680000 0.255000 1.010000 0.715000 ;
        RECT 0.680000 1.665000 1.010000 2.465000 ;
        RECT 1.520000 0.255000 1.850000 0.715000 ;
        RECT 1.520000 1.665000 1.850000 2.465000 ;
        RECT 2.360000 0.255000 2.690000 0.715000 ;
        RECT 2.360000 1.665000 2.690000 2.465000 ;
        RECT 3.200000 0.255000 3.530000 0.715000 ;
        RECT 3.200000 1.665000 3.530000 2.465000 ;
        RECT 3.735000 0.905000 4.055000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.255000  0.085000 0.510000 0.545000 ;
      RECT 0.255000  1.835000 0.510000 2.635000 ;
      RECT 1.180000  0.085000 1.350000 0.545000 ;
      RECT 1.180000  1.835000 1.350000 2.635000 ;
      RECT 2.020000  0.085000 2.190000 0.545000 ;
      RECT 2.020000  1.835000 2.190000 2.635000 ;
      RECT 2.860000  0.085000 3.030000 0.545000 ;
      RECT 2.860000  1.835000 3.030000 2.635000 ;
      RECT 3.700000  0.085000 4.005000 0.545000 ;
      RECT 3.700000  1.835000 4.000000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__inv_8
MACRO sky130_fd_sc_hd__inv_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_12 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.970000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.680000 1.075000 5.270000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.673000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 5.895000 0.905000 ;
        RECT 0.085000 0.905000 0.510000 1.495000 ;
        RECT 0.085000 1.495000 5.895000 1.665000 ;
        RECT 0.680000 0.255000 1.010000 0.715000 ;
        RECT 0.680000 1.665000 1.010000 2.465000 ;
        RECT 1.520000 0.255000 1.850000 0.715000 ;
        RECT 1.520000 1.665000 1.850000 2.465000 ;
        RECT 2.360000 0.255000 2.690000 0.715000 ;
        RECT 2.360000 1.665000 2.690000 2.465000 ;
        RECT 3.200000 0.255000 3.530000 0.715000 ;
        RECT 3.200000 1.665000 3.530000 2.465000 ;
        RECT 4.040000 0.255000 4.370000 0.715000 ;
        RECT 4.040000 1.665000 4.370000 2.465000 ;
        RECT 4.880000 0.255000 5.210000 0.715000 ;
        RECT 4.880000 1.665000 5.210000 2.465000 ;
        RECT 5.545000 0.905000 5.895000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.255000  0.085000 0.510000 0.545000 ;
      RECT 0.255000  1.835000 0.510000 2.635000 ;
      RECT 1.180000  0.085000 1.350000 0.545000 ;
      RECT 1.180000  1.835000 1.350000 2.635000 ;
      RECT 2.020000  0.085000 2.190000 0.545000 ;
      RECT 2.020000  1.835000 2.190000 2.635000 ;
      RECT 2.860000  0.085000 3.030000 0.545000 ;
      RECT 2.860000  1.835000 3.030000 2.635000 ;
      RECT 3.700000  0.085000 3.870000 0.545000 ;
      RECT 3.700000  1.835000 3.870000 2.635000 ;
      RECT 4.540000  0.085000 4.710000 0.545000 ;
      RECT 4.540000  1.835000 4.710000 2.635000 ;
      RECT 5.555000  0.085000 5.895000 0.545000 ;
      RECT 5.555000  1.835000 5.895000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__inv_12
MACRO sky130_fd_sc_hd__inv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  3.960000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 5.525000 1.315000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.580000 0.255000 0.910000 0.715000 ;
        RECT 0.580000 0.715000 6.790000 0.905000 ;
        RECT 0.580000 1.495000 6.790000 1.665000 ;
        RECT 0.580000 1.665000 0.910000 2.465000 ;
        RECT 1.420000 0.255000 1.750000 0.715000 ;
        RECT 1.420000 1.665000 1.750000 2.465000 ;
        RECT 2.260000 0.255000 2.590000 0.715000 ;
        RECT 2.260000 1.665000 2.590000 2.465000 ;
        RECT 3.100000 0.255000 3.430000 0.715000 ;
        RECT 3.100000 1.665000 3.430000 2.465000 ;
        RECT 3.940000 0.255000 4.270000 0.715000 ;
        RECT 3.940000 1.665000 4.270000 2.465000 ;
        RECT 4.780000 0.255000 5.110000 0.715000 ;
        RECT 4.780000 1.665000 5.110000 2.465000 ;
        RECT 5.620000 0.255000 5.950000 0.715000 ;
        RECT 5.620000 1.665000 5.950000 2.465000 ;
        RECT 6.460000 0.255000 6.790000 0.715000 ;
        RECT 6.460000 0.905000 6.790000 1.495000 ;
        RECT 6.460000 1.665000 6.790000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.180000  0.085000 0.410000 0.885000 ;
      RECT 0.200000  1.485000 0.410000 2.635000 ;
      RECT 1.080000  0.085000 1.250000 0.545000 ;
      RECT 1.080000  1.835000 1.250000 2.635000 ;
      RECT 1.920000  0.085000 2.090000 0.545000 ;
      RECT 1.920000  1.835000 2.090000 2.635000 ;
      RECT 2.760000  0.085000 2.930000 0.545000 ;
      RECT 2.760000  1.835000 2.930000 2.635000 ;
      RECT 3.600000  0.085000 3.770000 0.545000 ;
      RECT 3.600000  1.835000 3.770000 2.635000 ;
      RECT 4.440000  0.085000 4.610000 0.545000 ;
      RECT 4.440000  1.835000 4.610000 2.635000 ;
      RECT 5.280000  0.085000 5.450000 0.545000 ;
      RECT 5.280000  1.835000 5.450000 2.635000 ;
      RECT 6.120000  0.085000 6.290000 0.545000 ;
      RECT 6.120000  1.835000 6.290000 2.635000 ;
      RECT 6.960000  0.085000 7.170000 0.885000 ;
      RECT 6.960000  1.835000 7.170000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__inv_16
MACRO sky130_fd_sc_hd__lpflow_bleeder_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_bleeder_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN SHORT
    ANTENNAGATEAREA  0.270000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.275000 1.040000 1.975000 1.730000 ;
    END
  END SHORT
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.285000  0.085000 0.615000 0.870000 ;
      RECT 2.145000  0.540000 2.475000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_bleeder_1
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.196500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.985000 1.275000 1.355000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.345000 0.760000 ;
        RECT 0.085000 0.760000 0.255000 1.560000 ;
        RECT 0.085000 1.560000 0.355000 2.465000 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.875000 0.855000 2.465000 ;
      LAYER mcon ;
        RECT 0.610000 2.125000 0.780000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 1.310000 2.340000 ;
        RECT 0.550000 2.080000 0.840000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.425000  1.060000 0.710000 1.390000 ;
      RECT 0.525000  0.085000 0.855000 0.465000 ;
      RECT 0.540000  0.635000 1.205000 0.805000 ;
      RECT 0.540000  0.805000 0.710000 1.060000 ;
      RECT 0.540000  1.390000 0.710000 1.535000 ;
      RECT 0.540000  1.535000 1.205000 1.705000 ;
      RECT 1.035000  0.255000 1.205000 0.635000 ;
      RECT 1.035000  1.705000 1.205000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_1
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.745000 0.785000 1.240000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.383400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.040000 0.255000 1.245000 0.655000 ;
        RECT 1.040000 0.655000 1.725000 0.825000 ;
        RECT 1.060000 1.750000 1.725000 1.970000 ;
        RECT 1.060000 1.970000 1.245000 2.435000 ;
        RECT 1.385000 0.825000 1.725000 1.750000 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.855000 0.855000 2.465000 ;
      LAYER mcon ;
        RECT 0.610000 2.125000 0.780000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.415000 2.140000 1.750000 2.465000 ;
      LAYER mcon ;
        RECT 1.495000 2.140000 1.665000 2.310000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 1.770000 2.340000 ;
        RECT 0.550000 2.080000 0.840000 2.140000 ;
        RECT 1.435000 2.080000 1.725000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.585000 ;
      RECT 0.085000  0.585000 0.255000 1.410000 ;
      RECT 0.085000  1.410000 1.215000 1.580000 ;
      RECT 0.085000  1.580000 0.355000 2.435000 ;
      RECT 0.555000  0.085000 0.830000 0.565000 ;
      RECT 0.965000  0.995000 1.215000 1.410000 ;
      RECT 1.415000  0.085000 1.750000 0.485000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_2
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.755000 0.775000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.795200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.345000 1.305000 0.735000 ;
        RECT 1.010000 0.735000 2.660000 0.905000 ;
        RECT 1.025000 1.835000 2.165000 1.965000 ;
        RECT 1.025000 1.965000 1.390000 1.970000 ;
        RECT 1.025000 1.970000 1.385000 1.975000 ;
        RECT 1.025000 1.975000 1.370000 1.980000 ;
        RECT 1.025000 1.980000 1.330000 2.000000 ;
        RECT 1.025000 2.000000 1.325000 2.005000 ;
        RECT 1.025000 2.005000 1.265000 2.465000 ;
        RECT 1.185000 1.825000 2.165000 1.835000 ;
        RECT 1.195000 1.820000 2.165000 1.825000 ;
        RECT 1.205000 1.815000 2.165000 1.820000 ;
        RECT 1.215000 1.805000 2.165000 1.815000 ;
        RECT 1.245000 1.785000 2.165000 1.805000 ;
        RECT 1.270000 1.750000 2.165000 1.785000 ;
        RECT 1.905000 0.345000 2.165000 0.735000 ;
        RECT 1.905000 1.415000 2.660000 1.585000 ;
        RECT 1.905000 1.585000 2.165000 1.750000 ;
        RECT 1.935000 1.965000 2.165000 2.465000 ;
        RECT 2.255000 0.905000 2.660000 1.415000 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.835000 0.855000 2.465000 ;
      LAYER mcon ;
        RECT 0.610000 2.125000 0.780000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.435000 2.140000 1.765000 2.465000 ;
        RECT 2.335000 1.765000 2.620000 2.465000 ;
      LAYER mcon ;
        RECT 1.495000 2.140000 1.665000 2.310000 ;
        RECT 2.375000 2.125000 2.545000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 2.690000 2.340000 ;
        RECT 0.550000 2.080000 0.840000 2.140000 ;
        RECT 1.435000 2.080000 1.725000 2.140000 ;
        RECT 2.315000 2.080000 2.605000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.255000 0.385000 0.585000 ;
      RECT 0.085000  0.585000 0.255000 1.495000 ;
      RECT 0.085000  1.495000 1.115000 1.665000 ;
      RECT 0.085000  1.665000 0.355000 2.465000 ;
      RECT 0.555000  0.085000 0.830000 0.565000 ;
      RECT 0.945000  1.075000 2.085000 1.245000 ;
      RECT 0.945000  1.245000 1.115000 1.495000 ;
      RECT 1.475000  0.085000 1.730000 0.565000 ;
      RECT 2.335000  0.085000 2.615000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_4
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.426000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 0.400000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.590400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.420000 0.280000 1.680000 0.735000 ;
        RECT 1.420000 0.735000 4.730000 0.905000 ;
        RECT 1.420000 1.495000 4.730000 1.735000 ;
        RECT 1.420000 1.735000 1.680000 2.460000 ;
        RECT 2.280000 0.280000 2.540000 0.735000 ;
        RECT 2.280000 1.735000 2.540000 2.460000 ;
        RECT 3.140000 0.280000 3.400000 0.735000 ;
        RECT 3.140000 1.735000 3.400000 2.460000 ;
        RECT 3.760000 0.905000 4.730000 1.495000 ;
        RECT 4.000000 0.280000 4.260000 0.735000 ;
        RECT 4.000000 1.735000 4.260000 2.460000 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.525000 0.390000 2.465000 ;
      LAYER mcon ;
        RECT 0.175000 2.125000 0.345000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.990000 1.525000 1.250000 2.465000 ;
      LAYER mcon ;
        RECT 1.035000 2.125000 1.205000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.850000 1.905000 2.110000 2.465000 ;
      LAYER mcon ;
        RECT 1.890000 2.125000 2.060000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.710000 1.905000 2.970000 2.465000 ;
      LAYER mcon ;
        RECT 2.740000 2.125000 2.910000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.570000 1.905000 3.830000 2.465000 ;
      LAYER mcon ;
        RECT 3.620000 2.125000 3.790000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.430000 1.905000 4.725000 2.465000 ;
      LAYER mcon ;
        RECT 4.480000 2.125000 4.650000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 4.990000 2.340000 ;
        RECT 0.115000 2.080000 0.405000 2.140000 ;
        RECT 0.975000 2.080000 1.265000 2.140000 ;
        RECT 1.830000 2.080000 2.120000 2.140000 ;
        RECT 2.680000 2.080000 2.970000 2.140000 ;
        RECT 3.560000 2.080000 3.850000 2.140000 ;
        RECT 4.420000 2.080000 4.710000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.145000  0.085000 0.390000 0.545000 ;
      RECT 0.570000  0.265000 0.820000 1.075000 ;
      RECT 0.570000  1.075000 3.590000 1.325000 ;
      RECT 0.570000  1.325000 0.820000 2.460000 ;
      RECT 0.990000  0.085000 1.250000 0.610000 ;
      RECT 1.850000  0.085000 2.110000 0.565000 ;
      RECT 2.710000  0.085000 2.970000 0.565000 ;
      RECT 3.570000  0.085000 3.830000 0.565000 ;
      RECT 4.430000  0.085000 4.730000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_8
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.852000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.400000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.180800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.280000 0.280000 2.540000 0.735000 ;
        RECT 2.280000 0.735000 9.025000 0.905000 ;
        RECT 2.315000 1.495000 9.025000 1.720000 ;
        RECT 2.315000 1.720000 7.685000 1.735000 ;
        RECT 2.315000 1.735000 2.540000 2.460000 ;
        RECT 3.140000 0.280000 3.400000 0.735000 ;
        RECT 3.140000 1.735000 3.400000 2.460000 ;
        RECT 4.000000 0.280000 4.260000 0.735000 ;
        RECT 4.000000 1.735000 4.260000 2.460000 ;
        RECT 4.845000 0.280000 5.120000 0.735000 ;
        RECT 4.860000 1.735000 5.120000 2.460000 ;
        RECT 5.705000 0.280000 5.965000 0.735000 ;
        RECT 5.705000 1.735000 5.965000 2.460000 ;
        RECT 6.565000 0.280000 6.825000 0.735000 ;
        RECT 6.565000 1.735000 6.825000 2.460000 ;
        RECT 7.425000 0.280000 7.685000 0.735000 ;
        RECT 7.425000 1.735000 7.685000 2.460000 ;
        RECT 7.860000 0.905000 9.025000 1.495000 ;
        RECT 8.295000 0.280000 8.555000 0.735000 ;
        RECT 8.295000 1.720000 8.585000 2.460000 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.495000 0.425000 2.465000 ;
      LAYER mcon ;
        RECT 0.175000 2.125000 0.345000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.955000 1.495000 1.285000 2.465000 ;
      LAYER mcon ;
        RECT 1.035000 2.125000 1.205000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.815000 1.495000 2.145000 2.465000 ;
      LAYER mcon ;
        RECT 1.890000 2.125000 2.060000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.710000 1.905000 2.970000 2.465000 ;
      LAYER mcon ;
        RECT 2.740000 2.125000 2.910000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.570000 1.905000 3.830000 2.465000 ;
      LAYER mcon ;
        RECT 3.620000 2.125000 3.790000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.430000 1.905000 4.690000 2.465000 ;
      LAYER mcon ;
        RECT 4.480000 2.125000 4.650000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.290000 1.905000 5.535000 2.465000 ;
      LAYER mcon ;
        RECT 5.335000 2.125000 5.505000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.150000 1.905000 6.395000 2.465000 ;
      LAYER mcon ;
        RECT 6.195000 2.125000 6.365000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.010000 1.905000 7.255000 2.465000 ;
      LAYER mcon ;
        RECT 7.050000 2.125000 7.220000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.870000 1.905000 8.125000 2.465000 ;
      LAYER mcon ;
        RECT 7.900000 2.125000 8.070000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.755000 1.890000 9.025000 2.465000 ;
      LAYER mcon ;
        RECT 8.780000 2.125000 8.950000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 9.130000 2.340000 ;
        RECT 0.115000 2.080000 0.405000 2.140000 ;
        RECT 0.975000 2.080000 1.265000 2.140000 ;
        RECT 1.830000 2.080000 2.120000 2.140000 ;
        RECT 2.680000 2.080000 2.970000 2.140000 ;
        RECT 3.560000 2.080000 3.850000 2.140000 ;
        RECT 4.420000 2.080000 4.710000 2.140000 ;
        RECT 5.275000 2.080000 5.565000 2.140000 ;
        RECT 6.135000 2.080000 6.425000 2.140000 ;
        RECT 6.990000 2.080000 7.280000 2.140000 ;
        RECT 7.840000 2.080000 8.130000 2.140000 ;
        RECT 8.720000 2.080000 9.010000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.085000  0.085000 0.390000 0.595000 ;
      RECT 0.595000  0.265000 0.820000 1.075000 ;
      RECT 0.595000  1.075000 7.690000 1.325000 ;
      RECT 0.595000  1.325000 0.785000 2.465000 ;
      RECT 0.990000  0.085000 1.250000 0.610000 ;
      RECT 1.430000  0.265000 1.680000 1.075000 ;
      RECT 1.455000  1.325000 1.645000 2.460000 ;
      RECT 1.850000  0.085000 2.110000 0.645000 ;
      RECT 2.710000  0.085000 2.970000 0.565000 ;
      RECT 3.570000  0.085000 3.830000 0.565000 ;
      RECT 4.430000  0.085000 4.675000 0.565000 ;
      RECT 5.290000  0.085000 5.535000 0.565000 ;
      RECT 6.145000  0.085000 6.395000 0.565000 ;
      RECT 7.005000  0.085000 7.255000 0.565000 ;
      RECT 7.865000  0.085000 8.125000 0.565000 ;
      RECT 8.725000  0.085000 9.025000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_16
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.375000 0.325000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.336000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.590000 0.255000 0.840000 0.760000 ;
        RECT 0.590000 0.760000 1.295000 0.945000 ;
        RECT 0.595000 0.945000 1.295000 1.290000 ;
        RECT 0.595000 1.290000 0.765000 2.465000 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.665000 0.425000 2.465000 ;
      LAYER mcon ;
        RECT 0.155000 2.125000 0.325000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.935000 1.665000 1.295000 2.465000 ;
      LAYER mcon ;
        RECT 1.055000 2.125000 1.225000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 1.310000 2.340000 ;
        RECT 0.095000 2.080000 0.385000 2.140000 ;
        RECT 0.995000 2.080000 1.285000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 1.010000  0.085000 1.295000 0.590000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_1
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.576000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.065000 1.305000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.662600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.460000 1.755000 1.630000 ;
        RECT 0.155000 1.630000 0.375000 2.435000 ;
        RECT 1.025000 0.280000 1.250000 0.725000 ;
        RECT 1.025000 0.725000 1.755000 0.895000 ;
        RECT 1.045000 1.630000 1.235000 2.435000 ;
        RECT 1.475000 0.895000 1.755000 1.460000 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.800000 0.875000 2.465000 ;
      LAYER mcon ;
        RECT 0.600000 2.125000 0.770000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.405000 1.800000 1.735000 2.465000 ;
      LAYER mcon ;
        RECT 1.500000 2.125000 1.670000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 1.770000 2.340000 ;
        RECT 0.540000 2.080000 0.830000 2.140000 ;
        RECT 1.440000 2.080000 1.730000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.560000  0.085000 0.855000 0.610000 ;
      RECT 1.420000  0.085000 1.750000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_2
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.152000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.065000 2.660000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.075200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.725000 3.135000 0.895000 ;
        RECT 0.105000 0.895000 0.275000 1.460000 ;
        RECT 0.105000 1.460000 3.135000 1.630000 ;
        RECT 0.645000 1.630000 0.815000 2.435000 ;
        RECT 1.030000 0.280000 1.290000 0.725000 ;
        RECT 1.505000 1.630000 1.675000 2.435000 ;
        RECT 1.890000 0.280000 2.145000 0.725000 ;
        RECT 2.365000 1.630000 2.535000 2.435000 ;
        RECT 2.835000 0.895000 3.135000 1.460000 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.135000 1.800000 0.465000 2.465000 ;
      LAYER mcon ;
        RECT 0.195000 2.125000 0.365000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.995000 1.800000 1.325000 2.465000 ;
      LAYER mcon ;
        RECT 1.055000 2.125000 1.225000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.855000 1.800000 2.185000 2.465000 ;
      LAYER mcon ;
        RECT 1.955000 2.125000 2.125000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.715000 1.800000 3.045000 2.465000 ;
      LAYER mcon ;
        RECT 2.835000 2.125000 3.005000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 3.150000 2.340000 ;
        RECT 0.135000 2.080000 0.425000 2.140000 ;
        RECT 0.995000 2.080000 1.285000 2.140000 ;
        RECT 1.895000 2.080000 2.185000 2.140000 ;
        RECT 2.775000 2.080000 3.065000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.565000  0.085000 0.860000 0.555000 ;
      RECT 1.460000  0.085000 1.720000 0.555000 ;
      RECT 2.315000  0.085000 2.615000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_4
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.304000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.035000 4.865000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.090400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.695000 5.440000 0.865000 ;
        RECT 0.115000 0.865000 0.285000 1.460000 ;
        RECT 0.115000 1.460000 5.440000 1.630000 ;
        RECT 0.595000 1.630000 0.765000 2.435000 ;
        RECT 1.440000 1.630000 1.610000 2.435000 ;
        RECT 1.535000 0.280000 1.725000 0.695000 ;
        RECT 2.280000 1.630000 2.450000 2.435000 ;
        RECT 2.395000 0.280000 2.585000 0.695000 ;
        RECT 3.120000 1.630000 3.290000 2.435000 ;
        RECT 3.255000 0.280000 3.445000 0.695000 ;
        RECT 3.960000 1.630000 4.130000 2.435000 ;
        RECT 4.115000 0.280000 4.305000 0.695000 ;
        RECT 4.800000 1.630000 4.970000 2.435000 ;
        RECT 5.170000 0.865000 5.440000 1.460000 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.800000 0.425000 2.465000 ;
        RECT 5.140000 1.800000 5.470000 2.465000 ;
      LAYER mcon ;
        RECT 0.130000 2.125000 0.300000 2.295000 ;
        RECT 5.255000 2.125000 5.425000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.940000 1.800000 1.270000 2.465000 ;
      LAYER mcon ;
        RECT 0.990000 2.125000 1.160000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.780000 1.800000 2.110000 2.465000 ;
      LAYER mcon ;
        RECT 1.890000 2.125000 2.060000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.620000 1.800000 2.950000 2.465000 ;
      LAYER mcon ;
        RECT 2.770000 2.125000 2.940000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.460000 1.800000 3.790000 2.465000 ;
      LAYER mcon ;
        RECT 3.495000 2.125000 3.665000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.300000 1.800000 4.630000 2.465000 ;
      LAYER mcon ;
        RECT 4.355000 2.125000 4.525000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.080000 0.360000 2.140000 ;
        RECT 0.070000 2.140000 5.910000 2.340000 ;
        RECT 0.930000 2.080000 1.220000 2.140000 ;
        RECT 1.830000 2.080000 2.120000 2.140000 ;
        RECT 2.710000 2.080000 3.000000 2.140000 ;
        RECT 3.435000 2.080000 3.725000 2.140000 ;
        RECT 4.295000 2.080000 4.585000 2.140000 ;
        RECT 5.195000 2.080000 5.485000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 1.035000  0.085000 1.365000 0.525000 ;
      RECT 1.895000  0.085000 2.225000 0.525000 ;
      RECT 2.755000  0.085000 3.085000 0.525000 ;
      RECT 3.615000  0.085000 3.945000 0.525000 ;
      RECT 4.475000  0.085000 4.805000 0.525000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_8
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  4.608000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.345000 0.895000  2.155000 1.275000 ;
        RECT 8.930000 0.895000 10.710000 1.275000 ;
      LAYER mcon ;
        RECT 1.525000 1.105000 1.695000 1.275000 ;
        RECT 1.985000 1.105000 2.155000 1.275000 ;
        RECT 9.345000 1.105000 9.515000 1.275000 ;
        RECT 9.805000 1.105000 9.975000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465000 1.075000  2.215000 1.120000 ;
        RECT 1.465000 1.120000 10.035000 1.260000 ;
        RECT 1.465000 1.260000  2.215000 1.305000 ;
        RECT 9.285000 1.075000 10.035000 1.120000 ;
        RECT 9.285000 1.260000 10.035000 1.305000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  4.520900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.615000 1.455000 10.480000 1.665000 ;
        RECT  0.615000 1.665000  0.785000 2.465000 ;
        RECT  1.475000 1.665000  1.645000 2.465000 ;
        RECT  2.325000 0.280000  2.550000 1.415000 ;
        RECT  2.325000 1.415000  8.755000 1.455000 ;
        RECT  2.335000 1.665000  2.505000 2.465000 ;
        RECT  3.155000 0.280000  3.410000 1.415000 ;
        RECT  3.195000 1.665000  3.365000 2.465000 ;
        RECT  4.015000 0.280000  4.255000 1.415000 ;
        RECT  4.055000 1.665000  4.225000 2.465000 ;
        RECT  4.905000 0.280000  5.255000 1.415000 ;
        RECT  5.080000 1.665000  5.250000 2.465000 ;
        RECT  5.925000 0.280000  6.175000 1.415000 ;
        RECT  5.965000 1.665000  6.135000 2.465000 ;
        RECT  6.785000 0.280000  7.035000 1.415000 ;
        RECT  6.825000 1.665000  6.995000 2.465000 ;
        RECT  7.645000 0.280000  7.895000 1.415000 ;
        RECT  7.685000 1.665000  7.855000 2.465000 ;
        RECT  8.505000 0.280000  8.755000 1.415000 ;
        RECT  8.545000 1.665000  8.715000 2.465000 ;
        RECT  9.405000 1.665000  9.575000 2.465000 ;
        RECT 10.265000 1.665000 10.435000 2.465000 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.110000 1.495000  0.440000 2.465000 ;
        RECT 10.610000 1.835000 10.940000 2.465000 ;
      LAYER mcon ;
        RECT  0.130000 2.125000  0.300000 2.295000 ;
        RECT 10.720000 2.125000 10.890000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.965000 1.835000 1.295000 2.465000 ;
      LAYER mcon ;
        RECT 0.990000 2.125000 1.160000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.825000 1.835000 2.155000 2.465000 ;
      LAYER mcon ;
        RECT 1.890000 2.125000 2.060000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.685000 1.835000 3.015000 2.465000 ;
      LAYER mcon ;
        RECT 2.770000 2.125000 2.940000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.545000 1.835000 3.875000 2.465000 ;
      LAYER mcon ;
        RECT 3.690000 2.125000 3.860000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.425000 1.835000 4.755000 2.465000 ;
      LAYER mcon ;
        RECT 4.550000 2.125000 4.720000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.450000 1.835000 5.780000 2.465000 ;
      LAYER mcon ;
        RECT 5.450000 2.125000 5.620000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.315000 1.835000 6.645000 2.465000 ;
      LAYER mcon ;
        RECT 6.370000 2.125000 6.540000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.175000 1.835000 7.505000 2.465000 ;
      LAYER mcon ;
        RECT 7.230000 2.125000 7.400000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.035000 1.835000 8.365000 2.465000 ;
      LAYER mcon ;
        RECT 8.130000 2.125000 8.300000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.895000 1.835000 9.225000 2.465000 ;
      LAYER mcon ;
        RECT 8.960000 2.125000 9.130000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755000 1.835000 10.085000 2.465000 ;
      LAYER mcon ;
        RECT 9.820000 2.125000 9.990000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT  0.070000 2.080000  0.360000 2.140000 ;
        RECT  0.070000 2.140000 10.970000 2.340000 ;
        RECT  0.930000 2.080000  1.220000 2.140000 ;
        RECT  1.830000 2.080000  2.120000 2.140000 ;
        RECT  2.710000 2.080000  3.000000 2.140000 ;
        RECT  3.630000 2.080000  3.920000 2.140000 ;
        RECT  4.490000 2.080000  4.780000 2.140000 ;
        RECT  5.390000 2.080000  5.680000 2.140000 ;
        RECT  6.310000 2.080000  6.600000 2.140000 ;
        RECT  7.170000 2.080000  7.460000 2.140000 ;
        RECT  8.070000 2.080000  8.360000 2.140000 ;
        RECT  8.900000 2.080000  9.190000 2.140000 ;
        RECT  9.760000 2.080000 10.050000 2.140000 ;
        RECT 10.660000 2.080000 10.950000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 11.040000 0.085000 ;
      RECT 0.000000  2.635000 11.040000 2.805000 ;
      RECT 1.855000  0.085000  2.125000 0.610000 ;
      RECT 2.720000  0.085000  2.985000 0.610000 ;
      RECT 3.580000  0.085000  3.845000 0.610000 ;
      RECT 4.465000  0.085000  4.730000 0.610000 ;
      RECT 5.490000  0.085000  5.755000 0.610000 ;
      RECT 6.350000  0.085000  6.575000 0.610000 ;
      RECT 7.210000  0.085000  7.475000 0.610000 ;
      RECT 8.070000  0.085000  8.335000 0.610000 ;
      RECT 8.930000  0.085000  9.195000 0.610000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_16
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_3
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_3 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.545000 1.295000 2.465000 ;
        RECT 0.775000 1.005000 1.295000 1.545000 ;
      LAYER mcon ;
        RECT 0.145000 2.125000 0.315000 2.295000 ;
        RECT 0.605000 2.125000 0.775000 2.295000 ;
        RECT 1.065000 2.125000 1.235000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 1.310000 2.340000 ;
        RECT 0.085000 2.080000 1.295000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.085000  0.085000 1.295000 0.835000 ;
      RECT 0.085000  0.835000 0.605000 1.375000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_3
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.545000 1.755000 2.465000 ;
        RECT 1.005000 1.025000 1.755000 1.545000 ;
      LAYER mcon ;
        RECT 0.145000 2.125000 0.315000 2.295000 ;
        RECT 0.605000 2.125000 0.775000 2.295000 ;
        RECT 1.065000 2.125000 1.235000 2.295000 ;
        RECT 1.525000 2.125000 1.695000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 1.770000 2.340000 ;
        RECT 0.085000 2.080000 1.755000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.085000  0.085000 1.755000 0.855000 ;
      RECT 0.085000  0.855000 0.835000 1.375000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_4
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_6 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.545000 2.675000 2.465000 ;
        RECT 1.465000 1.025000 2.675000 1.545000 ;
      LAYER mcon ;
        RECT 0.145000 2.125000 0.315000 2.295000 ;
        RECT 0.605000 2.125000 0.775000 2.295000 ;
        RECT 1.065000 2.125000 1.235000 2.295000 ;
        RECT 1.525000 2.125000 1.695000 2.295000 ;
        RECT 1.985000 2.125000 2.155000 2.295000 ;
        RECT 2.445000 2.125000 2.615000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 2.690000 2.340000 ;
        RECT 0.085000 2.080000 2.675000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.085000 2.675000 0.855000 ;
      RECT 0.085000  0.855000 1.295000 1.375000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_6
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.545000 3.595000 2.465000 ;
        RECT 1.905000 1.025000 3.595000 1.545000 ;
      LAYER mcon ;
        RECT 0.145000 2.125000 0.315000 2.295000 ;
        RECT 0.605000 2.125000 0.775000 2.295000 ;
        RECT 1.065000 2.125000 1.235000 2.295000 ;
        RECT 1.525000 2.125000 1.695000 2.295000 ;
        RECT 1.985000 2.125000 2.155000 2.295000 ;
        RECT 2.445000 2.125000 2.615000 2.295000 ;
        RECT 2.905000 2.125000 3.075000 2.295000 ;
        RECT 3.365000 2.125000 3.535000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 3.610000 2.340000 ;
        RECT 0.085000 2.080000 3.595000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.085000 3.595000 0.855000 ;
      RECT 0.085000  0.855000 1.735000 1.375000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_8
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_12 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.545000 5.430000 2.465000 ;
        RECT 2.835000 1.025000 5.430000 1.545000 ;
      LAYER mcon ;
        RECT 0.145000 2.125000 0.315000 2.295000 ;
        RECT 0.605000 2.125000 0.775000 2.295000 ;
        RECT 1.065000 2.125000 1.235000 2.295000 ;
        RECT 1.525000 2.125000 1.695000 2.295000 ;
        RECT 1.985000 2.125000 2.155000 2.295000 ;
        RECT 2.445000 2.125000 2.615000 2.295000 ;
        RECT 2.905000 2.125000 3.075000 2.295000 ;
        RECT 3.365000 2.125000 3.535000 2.295000 ;
        RECT 3.825000 2.125000 3.995000 2.295000 ;
        RECT 4.285000 2.125000 4.455000 2.295000 ;
        RECT 4.745000 2.125000 4.915000 2.295000 ;
        RECT 5.205000 2.125000 5.375000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 5.450000 2.340000 ;
        RECT 0.085000 2.080000 5.435000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.085000 5.430000 0.855000 ;
      RECT 0.085000  0.855000 2.665000 1.375000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_12
MACRO sky130_fd_sc_hd__lpflow_inputiso0n_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso0n_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.075000 0.775000 1.325000 ;
        RECT 0.100000 1.325000 0.365000 1.685000 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 1.075000 1.335000 1.325000 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  0.657000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655000 0.255000 2.215000 0.545000 ;
        RECT 1.755000 1.915000 2.215000 2.465000 ;
        RECT 1.965000 0.545000 2.215000 1.915000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.285000  0.355000 0.615000 0.715000 ;
      RECT 0.285000  0.715000 1.675000 0.905000 ;
      RECT 0.285000  1.965000 0.565000 2.635000 ;
      RECT 0.735000  1.575000 1.675000 1.745000 ;
      RECT 0.735000  1.745000 1.035000 2.295000 ;
      RECT 1.235000  0.085000 1.485000 0.545000 ;
      RECT 1.235000  1.915000 1.565000 2.635000 ;
      RECT 1.505000  0.905000 1.675000 0.995000 ;
      RECT 1.505000  0.995000 1.795000 1.325000 ;
      RECT 1.505000  1.325000 1.675000 1.575000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso0n_1
MACRO sky130_fd_sc_hd__lpflow_inputiso0p_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso0p_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 1.645000 2.175000 1.955000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.765000 0.445000 1.615000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.350000 1.580000 2.655000 2.365000 ;
        RECT 2.415000 0.255000 2.655000 0.775000 ;
        RECT 2.480000 0.775000 2.655000 1.580000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.590000 ;
      RECT 0.175000  1.785000 0.850000 2.015000 ;
      RECT 0.175000  2.015000 0.345000 2.445000 ;
      RECT 0.515000  2.185000 0.845000 2.635000 ;
      RECT 0.595000  0.280000 0.835000 0.655000 ;
      RECT 0.615000  0.655000 0.835000 0.805000 ;
      RECT 0.615000  0.805000 1.150000 1.135000 ;
      RECT 0.615000  1.135000 0.850000 1.785000 ;
      RECT 1.020000  1.305000 2.305000 1.325000 ;
      RECT 1.020000  1.325000 1.880000 1.475000 ;
      RECT 1.020000  1.475000 1.305000 2.420000 ;
      RECT 1.115000  0.270000 1.285000 0.415000 ;
      RECT 1.115000  0.415000 1.490000 0.610000 ;
      RECT 1.320000  0.610000 1.490000 0.945000 ;
      RECT 1.320000  0.945000 2.305000 1.305000 ;
      RECT 1.485000  2.165000 2.170000 2.635000 ;
      RECT 1.850000  0.085000 2.245000 0.580000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso0p_1
MACRO sky130_fd_sc_hd__lpflow_inputiso1n_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso1n_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 2.085000 1.735000 2.415000 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.425000 1.325000 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 0.415000 2.675000 0.760000 ;
        RECT 2.405000 1.495000 2.675000 2.465000 ;
        RECT 2.505000 0.760000 2.675000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.110000  0.265000 0.420000 0.735000 ;
      RECT 0.110000  0.735000 0.845000 0.905000 ;
      RECT 0.590000  0.085000 1.325000 0.565000 ;
      RECT 0.595000  0.905000 0.845000 0.995000 ;
      RECT 0.595000  0.995000 1.335000 1.325000 ;
      RECT 0.595000  1.325000 0.765000 1.885000 ;
      RECT 0.990000  1.495000 2.235000 1.665000 ;
      RECT 0.990000  1.665000 1.410000 1.915000 ;
      RECT 1.495000  0.305000 1.665000 0.655000 ;
      RECT 1.495000  0.655000 2.235000 0.825000 ;
      RECT 1.835000  0.085000 2.215000 0.485000 ;
      RECT 1.915000  1.835000 2.195000 2.635000 ;
      RECT 2.065000  0.825000 2.235000 0.995000 ;
      RECT 2.065000  0.995000 2.295000 1.325000 ;
      RECT 2.065000  1.325000 2.235000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso1n_1
MACRO sky130_fd_sc_hd__lpflow_inputiso1p_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso1p_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.765000 0.500000 1.325000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.765000 1.275000 1.325000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.509000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.255000 2.180000 0.825000 ;
        RECT 1.645000 1.845000 2.180000 2.465000 ;
        RECT 1.865000 0.825000 2.180000 1.845000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.250000  0.085000 0.490000 0.595000 ;
      RECT 0.270000  1.495000 1.695000 1.665000 ;
      RECT 0.270000  1.665000 0.660000 1.840000 ;
      RECT 0.670000  0.265000 0.950000 0.595000 ;
      RECT 0.670000  0.595000 0.840000 1.495000 ;
      RECT 1.145000  1.835000 1.475000 2.635000 ;
      RECT 1.180000  0.085000 1.395000 0.595000 ;
      RECT 1.525000  0.995000 1.695000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso1p_1
MACRO sky130_fd_sc_hd__lpflow_inputisolatch_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputisolatch_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.750000 0.765000 2.125000 1.095000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.690000 0.415000 4.975000 0.745000 ;
        RECT 4.690000 1.670000 4.975000 2.455000 ;
        RECT 4.805000 0.745000 4.975000 1.670000 ;
    END
  END Q
  PIN SLEEP_B
    ANTENNAGATEAREA  0.145500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.985000 0.330000 1.625000 ;
    END
  END SLEEP_B
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.130000 ;
      RECT 0.610000  1.130000 0.810000 1.460000 ;
      RECT 0.610000  1.460000 0.780000 1.795000 ;
      RECT 0.980000  0.740000 1.185000 0.910000 ;
      RECT 0.980000  0.910000 1.150000 1.825000 ;
      RECT 0.980000  1.825000 1.185000 1.915000 ;
      RECT 0.980000  1.915000 2.845000 1.965000 ;
      RECT 1.015000  0.345000 1.185000 0.740000 ;
      RECT 1.015000  1.965000 2.845000 2.085000 ;
      RECT 1.015000  2.085000 1.185000 2.465000 ;
      RECT 1.320000  1.240000 1.490000 1.525000 ;
      RECT 1.320000  1.525000 2.335000 1.695000 ;
      RECT 1.455000  0.085000 1.785000 0.465000 ;
      RECT 1.455000  2.255000 1.850000 2.635000 ;
      RECT 2.050000  1.355000 2.335000 1.525000 ;
      RECT 2.295000  0.705000 2.675000 1.035000 ;
      RECT 2.310000  2.255000 3.185000 2.425000 ;
      RECT 2.380000  0.365000 3.040000 0.535000 ;
      RECT 2.505000  1.035000 2.675000 1.575000 ;
      RECT 2.505000  1.575000 2.845000 1.915000 ;
      RECT 2.870000  0.535000 3.040000 0.995000 ;
      RECT 2.870000  0.995000 3.780000 1.165000 ;
      RECT 3.015000  1.165000 3.780000 1.325000 ;
      RECT 3.015000  1.325000 3.185000 2.255000 ;
      RECT 3.265000  0.085000 3.595000 0.530000 ;
      RECT 3.355000  2.135000 3.525000 2.635000 ;
      RECT 3.420000  1.535000 4.125000 1.865000 ;
      RECT 3.835000  0.415000 4.125000 0.745000 ;
      RECT 3.835000  1.865000 4.125000 2.435000 ;
      RECT 3.950000  0.745000 4.125000 1.535000 ;
      RECT 4.295000  0.085000 4.465000 0.715000 ;
      RECT 4.295000  1.570000 4.465000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_inputisolatch_1
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.725000 0.325000 1.325000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.960000 1.065000 1.325000 1.325000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.235000 0.255000 1.565000 0.725000 ;
        RECT 1.235000 0.725000 2.215000 0.895000 ;
        RECT 1.655000 1.850000 2.215000 2.465000 ;
        RECT 2.035000 0.895000 2.215000 1.850000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.330000  0.370000 0.675000 0.545000 ;
      RECT 0.415000  1.510000 1.705000 1.680000 ;
      RECT 0.415000  1.680000 0.675000 1.905000 ;
      RECT 0.495000  0.545000 0.675000 1.510000 ;
      RECT 0.855000  0.085000 1.065000 0.895000 ;
      RECT 0.875000  1.855000 1.205000 2.635000 ;
      RECT 1.535000  1.075000 1.865000 1.245000 ;
      RECT 1.535000  1.245000 1.705000 1.510000 ;
      RECT 1.735000  0.085000 2.120000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_1
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.600000 1.065000 3.125000 1.275000 ;
        RECT 2.910000 1.275000 3.125000 1.965000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.480000 1.065000 0.920000 1.275000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 1.705000 0.895000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 1.415000 0.895000 1.665000 2.125000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.085000 0.365000 0.895000 ;
      RECT 0.085000  1.445000 1.245000 1.655000 ;
      RECT 0.085000  1.655000 0.405000 2.465000 ;
      RECT 0.575000  1.825000 0.825000 2.635000 ;
      RECT 0.995000  1.655000 1.245000 2.295000 ;
      RECT 0.995000  2.295000 2.125000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.835000  1.445000 2.090000 1.890000 ;
      RECT 1.835000  1.890000 2.125000 2.295000 ;
      RECT 1.875000  0.085000 2.045000 0.895000 ;
      RECT 1.875000  1.075000 2.430000 1.245000 ;
      RECT 2.215000  0.725000 2.565000 0.895000 ;
      RECT 2.215000  0.895000 2.430000 1.075000 ;
      RECT 2.260000  1.245000 2.430000 1.445000 ;
      RECT 2.260000  1.445000 2.565000 1.615000 ;
      RECT 2.395000  0.445000 2.565000 0.725000 ;
      RECT 2.395000  1.615000 2.565000 2.460000 ;
      RECT 2.775000  0.085000 3.030000 0.845000 ;
      RECT 2.775000  2.145000 3.025000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_2
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.075000 4.975000 1.320000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.360000 1.075000 1.800000 1.275000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 3.385000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.215000 0.255000 2.545000 0.725000 ;
        RECT 2.295000 0.905000 2.625000 1.445000 ;
        RECT 2.295000 1.445000 3.305000 1.745000 ;
        RECT 2.295000 1.745000 2.465000 2.125000 ;
        RECT 3.055000 0.255000 3.385000 0.725000 ;
        RECT 3.135000 1.745000 3.305000 2.125000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.085000 0.365000 0.905000 ;
      RECT 0.085000  1.455000 2.125000 1.665000 ;
      RECT 0.085000  1.665000 0.365000 2.465000 ;
      RECT 0.535000  1.835000 0.865000 2.635000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.035000  1.665000 1.205000 2.465000 ;
      RECT 1.375000  1.835000 1.625000 2.635000 ;
      RECT 1.795000  1.665000 2.125000 2.295000 ;
      RECT 1.795000  2.295000 3.855000 2.465000 ;
      RECT 1.875000  0.085000 2.045000 0.555000 ;
      RECT 2.635000  1.935000 2.965000 2.295000 ;
      RECT 2.715000  0.085000 2.885000 0.555000 ;
      RECT 2.795000  1.075000 4.275000 1.275000 ;
      RECT 3.475000  1.575000 3.855000 2.295000 ;
      RECT 3.555000  0.085000 3.845000 0.905000 ;
      RECT 4.025000  0.255000 4.355000 0.815000 ;
      RECT 4.025000  0.815000 4.275000 1.075000 ;
      RECT 4.025000  1.275000 4.275000 1.575000 ;
      RECT 4.025000  1.575000 4.355000 2.465000 ;
      RECT 4.525000  0.085000 4.815000 0.905000 ;
      RECT 4.525000  1.495000 4.930000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_4
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.265000 1.065000 ;
        RECT 0.085000 1.065000 0.575000 1.285000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.270000 1.075000 8.010000 1.275000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  2.484000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005000 0.255000 2.335000 0.725000 ;
        RECT 2.005000 0.725000 8.655000 0.905000 ;
        RECT 2.845000 0.255000 3.175000 0.725000 ;
        RECT 3.685000 0.255000 4.015000 0.725000 ;
        RECT 4.525000 0.255000 4.855000 0.725000 ;
        RECT 5.365000 0.255000 5.695000 0.725000 ;
        RECT 5.405000 1.445000 8.655000 1.615000 ;
        RECT 5.405000 1.615000 5.655000 2.125000 ;
        RECT 6.205000 0.255000 6.535000 0.725000 ;
        RECT 6.245000 1.615000 6.495000 2.125000 ;
        RECT 7.045000 0.255000 7.375000 0.725000 ;
        RECT 7.085000 1.615000 7.335000 2.125000 ;
        RECT 7.885000 0.255000 8.215000 0.725000 ;
        RECT 7.925000 1.615000 8.175000 2.125000 ;
        RECT 8.180000 0.905000 8.655000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.930000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.195000  1.455000 0.415000 2.635000 ;
      RECT 0.435000  0.085000 0.655000 0.895000 ;
      RECT 0.585000  1.455000 0.915000 2.465000 ;
      RECT 0.745000  1.065000 1.155000 1.075000 ;
      RECT 0.745000  1.075000 5.000000 1.285000 ;
      RECT 0.745000  1.285000 0.915000 1.455000 ;
      RECT 0.825000  0.255000 1.155000 1.065000 ;
      RECT 1.085000  1.455000 1.330000 2.635000 ;
      RECT 1.325000  0.085000 1.835000 0.905000 ;
      RECT 1.555000  1.455000 5.235000 1.665000 ;
      RECT 1.555000  1.665000 1.875000 2.465000 ;
      RECT 2.045000  1.835000 2.295000 2.635000 ;
      RECT 2.465000  1.665000 2.715000 2.465000 ;
      RECT 2.505000  0.085000 2.675000 0.555000 ;
      RECT 2.885000  1.835000 3.135000 2.635000 ;
      RECT 3.305000  1.665000 3.555000 2.465000 ;
      RECT 3.345000  0.085000 3.515000 0.555000 ;
      RECT 3.725000  1.835000 3.975000 2.635000 ;
      RECT 4.145000  1.665000 4.395000 2.465000 ;
      RECT 4.185000  0.085000 4.355000 0.555000 ;
      RECT 4.565000  1.835000 4.815000 2.635000 ;
      RECT 4.985000  1.665000 5.235000 2.295000 ;
      RECT 4.985000  2.295000 8.595000 2.465000 ;
      RECT 5.025000  0.085000 5.195000 0.555000 ;
      RECT 5.825000  1.785000 6.075000 2.295000 ;
      RECT 5.865000  0.085000 6.035000 0.555000 ;
      RECT 6.665000  1.785000 6.915000 2.295000 ;
      RECT 6.705000  0.085000 6.875000 0.555000 ;
      RECT 7.505000  1.785000 7.755000 2.295000 ;
      RECT 7.545000  0.085000 7.715000 0.555000 ;
      RECT 8.345000  1.785000 8.595000 2.295000 ;
      RECT 8.385000  0.085000 8.655000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_8
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.56000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.315000 0.995000 ;
        RECT 0.085000 0.995000 0.665000 1.325000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  3.960000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.450000 1.075000 15.650000 1.285000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  4.968000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  2.925000 0.255000  3.255000 0.725000 ;
        RECT  2.925000 0.725000 16.475000 0.905000 ;
        RECT  3.765000 0.255000  4.095000 0.725000 ;
        RECT  4.605000 0.255000  4.935000 0.725000 ;
        RECT  5.445000 0.255000  5.775000 0.725000 ;
        RECT  6.285000 0.255000  6.615000 0.725000 ;
        RECT  7.125000 0.255000  7.455000 0.725000 ;
        RECT  7.965000 0.255000  8.295000 0.725000 ;
        RECT  8.805000 0.255000  9.135000 0.725000 ;
        RECT  9.645000 0.255000  9.975000 0.725000 ;
        RECT  9.685000 1.455000 16.475000 1.625000 ;
        RECT  9.685000 1.625000  9.935000 2.125000 ;
        RECT 10.485000 0.255000 10.815000 0.725000 ;
        RECT 10.525000 1.625000 10.775000 2.125000 ;
        RECT 11.325000 0.255000 11.655000 0.725000 ;
        RECT 11.365000 1.625000 11.615000 2.125000 ;
        RECT 12.165000 0.255000 12.495000 0.725000 ;
        RECT 12.205000 1.625000 12.455000 2.125000 ;
        RECT 13.005000 0.255000 13.335000 0.725000 ;
        RECT 13.045000 1.625000 13.295000 2.125000 ;
        RECT 13.845000 0.255000 14.175000 0.725000 ;
        RECT 13.885000 1.625000 14.135000 2.125000 ;
        RECT 14.685000 0.255000 15.015000 0.725000 ;
        RECT 14.725000 1.625000 14.975000 2.125000 ;
        RECT 15.525000 0.255000 15.855000 0.725000 ;
        RECT 15.565000 1.625000 15.815000 2.125000 ;
        RECT 15.820000 0.905000 16.475000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 16.560000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 16.750000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 16.560000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 16.560000 0.085000 ;
      RECT  0.000000  2.635000 16.560000 2.805000 ;
      RECT  0.300000  1.495000  0.515000 2.635000 ;
      RECT  0.485000  0.085000  0.815000 0.825000 ;
      RECT  0.685000  1.495000  1.015000 2.465000 ;
      RECT  0.835000  1.065000  2.035000 1.075000 ;
      RECT  0.835000  1.075000  9.280000 1.285000 ;
      RECT  0.835000  1.285000  1.015000 1.495000 ;
      RECT  0.985000  0.255000  1.195000 1.065000 ;
      RECT  1.185000  1.455000  1.355000 2.635000 ;
      RECT  1.365000  0.085000  1.615000 0.895000 ;
      RECT  1.525000  1.285000  1.855000 2.465000 ;
      RECT  1.785000  0.255000  2.035000 1.065000 ;
      RECT  2.025000  1.455000  2.270000 2.635000 ;
      RECT  2.205000  0.085000  2.755000 0.905000 ;
      RECT  2.475000  1.455000  9.515000 1.665000 ;
      RECT  2.475000  1.665000  2.795000 2.465000 ;
      RECT  2.965000  1.835000  3.215000 2.635000 ;
      RECT  3.385000  1.665000  3.635000 2.465000 ;
      RECT  3.425000  0.085000  3.595000 0.555000 ;
      RECT  3.805000  1.835000  4.055000 2.635000 ;
      RECT  4.225000  1.665000  4.475000 2.465000 ;
      RECT  4.265000  0.085000  4.435000 0.555000 ;
      RECT  4.645000  1.835000  4.895000 2.635000 ;
      RECT  5.065000  1.665000  5.315000 2.465000 ;
      RECT  5.105000  0.085000  5.275000 0.555000 ;
      RECT  5.485000  1.835000  5.735000 2.635000 ;
      RECT  5.905000  1.665000  6.155000 2.465000 ;
      RECT  5.945000  0.085000  6.115000 0.555000 ;
      RECT  6.325000  1.835000  6.575000 2.635000 ;
      RECT  6.745000  1.665000  6.995000 2.465000 ;
      RECT  6.785000  0.085000  6.955000 0.555000 ;
      RECT  7.165000  1.835000  7.415000 2.635000 ;
      RECT  7.585000  1.665000  7.835000 2.465000 ;
      RECT  7.625000  0.085000  7.795000 0.555000 ;
      RECT  8.005000  1.835000  8.255000 2.635000 ;
      RECT  8.425000  1.665000  8.675000 2.465000 ;
      RECT  8.465000  0.085000  8.635000 0.555000 ;
      RECT  8.845000  1.835000  9.095000 2.635000 ;
      RECT  9.265000  1.665000  9.515000 2.295000 ;
      RECT  9.265000  2.295000 16.235000 2.465000 ;
      RECT  9.305000  0.085000  9.475000 0.555000 ;
      RECT 10.105000  1.795000 10.355000 2.295000 ;
      RECT 10.145000  0.085000 10.315000 0.555000 ;
      RECT 10.945000  1.795000 11.195000 2.295000 ;
      RECT 10.985000  0.085000 11.155000 0.555000 ;
      RECT 11.785000  1.795000 12.035000 2.295000 ;
      RECT 11.825000  0.085000 11.995000 0.555000 ;
      RECT 12.625000  1.795000 12.875000 2.295000 ;
      RECT 12.665000  0.085000 12.835000 0.555000 ;
      RECT 13.465000  1.795000 13.715000 2.295000 ;
      RECT 13.505000  0.085000 13.675000 0.555000 ;
      RECT 14.305000  1.795000 14.555000 2.295000 ;
      RECT 14.345000  0.085000 14.515000 0.555000 ;
      RECT 15.145000  1.795000 15.395000 2.295000 ;
      RECT 15.185000  0.085000 15.355000 0.555000 ;
      RECT 15.985000  1.795000 16.235000 2.295000 ;
      RECT 16.025000  0.085000 16.295000 0.555000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_16
MACRO sky130_fd_sc_hd__lpflow_isobufsrckapwr_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrckapwr_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.26000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.615000 1.320000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.260000 1.075000 4.700000 1.275000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  3.180800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  7.340000 0.280000  7.600000 0.735000 ;
        RECT  7.340000 0.735000 14.085000 0.905000 ;
        RECT  7.375000 1.495000 14.085000 1.720000 ;
        RECT  7.375000 1.720000 12.745000 1.735000 ;
        RECT  7.375000 1.735000  7.600000 2.460000 ;
        RECT  8.200000 0.280000  8.460000 0.735000 ;
        RECT  8.200000 1.735000  8.460000 2.460000 ;
        RECT  9.060000 0.280000  9.320000 0.735000 ;
        RECT  9.060000 1.735000  9.320000 2.460000 ;
        RECT  9.905000 0.280000 10.180000 0.735000 ;
        RECT  9.920000 1.735000 10.180000 2.460000 ;
        RECT 10.765000 0.280000 11.025000 0.735000 ;
        RECT 10.765000 1.735000 11.025000 2.460000 ;
        RECT 11.625000 0.280000 11.885000 0.735000 ;
        RECT 11.625000 1.735000 11.885000 2.460000 ;
        RECT 12.485000 0.280000 12.745000 0.735000 ;
        RECT 12.485000 1.735000 12.745000 2.460000 ;
        RECT 12.920000 0.905000 14.085000 1.495000 ;
        RECT 13.355000 0.280000 13.615000 0.735000 ;
        RECT 13.355000 1.720000 13.645000 2.460000 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 10.350000 1.905000 10.595000 2.465000 ;
      LAYER mcon ;
        RECT 10.395000 2.125000 10.565000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 11.210000 1.905000 11.455000 2.465000 ;
      LAYER mcon ;
        RECT 11.255000 2.125000 11.425000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 12.070000 1.905000 12.315000 2.465000 ;
      LAYER mcon ;
        RECT 12.110000 2.125000 12.280000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 12.930000 1.905000 13.185000 2.465000 ;
      LAYER mcon ;
        RECT 12.960000 2.125000 13.130000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 13.815000 1.890000 14.085000 2.465000 ;
      LAYER mcon ;
        RECT 13.840000 2.125000 14.010000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.155000 1.495000 5.485000 2.465000 ;
      LAYER mcon ;
        RECT 5.235000 2.125000 5.405000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.015000 1.495000 6.345000 2.465000 ;
      LAYER mcon ;
        RECT 6.095000 2.125000 6.265000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.875000 1.495000 7.205000 2.465000 ;
      LAYER mcon ;
        RECT 6.950000 2.125000 7.120000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.770000 1.905000 8.030000 2.465000 ;
      LAYER mcon ;
        RECT 7.800000 2.125000 7.970000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.630000 1.905000 8.890000 2.465000 ;
      LAYER mcon ;
        RECT 8.680000 2.125000 8.850000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.490000 1.905000 9.750000 2.465000 ;
      LAYER mcon ;
        RECT 9.540000 2.125000 9.710000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT  0.070000 2.140000 14.190000 2.340000 ;
        RECT  5.175000 2.080000  5.465000 2.140000 ;
        RECT  6.035000 2.080000  6.325000 2.140000 ;
        RECT  6.890000 2.080000  7.180000 2.140000 ;
        RECT  7.740000 2.080000  8.030000 2.140000 ;
        RECT  8.620000 2.080000  8.910000 2.140000 ;
        RECT  9.480000 2.080000  9.770000 2.140000 ;
        RECT 10.335000 2.080000 10.625000 2.140000 ;
        RECT 11.195000 2.080000 11.485000 2.140000 ;
        RECT 12.050000 2.080000 12.340000 2.140000 ;
        RECT 12.900000 2.080000 13.190000 2.140000 ;
        RECT 13.780000 2.080000 14.070000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.260000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
    PORT
      LAYER pwell ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 14.450000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.260000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.260000 0.085000 ;
      RECT  0.000000  2.635000 14.260000 2.805000 ;
      RECT  0.130000  1.495000  0.535000 2.635000 ;
      RECT  0.245000  0.085000  0.535000 0.905000 ;
      RECT  0.705000  0.255000  1.035000 0.815000 ;
      RECT  0.705000  1.575000  1.035000 2.465000 ;
      RECT  0.785000  0.815000  1.035000 1.075000 ;
      RECT  0.785000  1.075000  2.265000 1.275000 ;
      RECT  0.785000  1.275000  1.035000 1.575000 ;
      RECT  1.205000  1.575000  1.585000 2.295000 ;
      RECT  1.205000  2.295000  3.265000 2.465000 ;
      RECT  1.215000  0.085000  1.505000 0.905000 ;
      RECT  1.675000  0.255000  2.005000 0.725000 ;
      RECT  1.675000  0.725000  4.525000 0.905000 ;
      RECT  1.755000  1.445000  2.765000 1.745000 ;
      RECT  1.755000  1.745000  1.925000 2.125000 ;
      RECT  2.095000  1.935000  2.425000 2.295000 ;
      RECT  2.175000  0.085000  2.345000 0.555000 ;
      RECT  2.435000  0.905000  3.095000 0.965000 ;
      RECT  2.435000  0.965000  2.765000 1.445000 ;
      RECT  2.515000  0.255000  2.845000 0.725000 ;
      RECT  2.595000  1.745000  2.765000 2.125000 ;
      RECT  2.935000  1.455000  4.975000 1.665000 ;
      RECT  2.935000  1.665000  3.265000 2.295000 ;
      RECT  3.015000  0.085000  3.185000 0.555000 ;
      RECT  3.355000  0.255000  3.685000 0.725000 ;
      RECT  3.435000  1.835000  3.685000 2.635000 ;
      RECT  3.855000  0.085000  4.025000 0.555000 ;
      RECT  3.855000  1.665000  4.025000 2.465000 ;
      RECT  4.195000  0.255000  4.525000 0.725000 ;
      RECT  4.195000  1.835000  4.525000 2.635000 ;
      RECT  4.695000  0.085000  5.450000 0.565000 ;
      RECT  4.695000  0.565000  4.975000 0.905000 ;
      RECT  4.695000  1.665000  4.975000 2.465000 ;
      RECT  5.145000  0.735000  5.460000 1.325000 ;
      RECT  5.655000  0.265000  5.880000 1.075000 ;
      RECT  5.655000  1.075000 12.750000 1.325000 ;
      RECT  5.655000  1.325000  5.845000 2.465000 ;
      RECT  6.050000  0.085000  6.310000 0.610000 ;
      RECT  6.490000  0.265000  6.740000 1.075000 ;
      RECT  6.515000  1.325000  6.705000 2.460000 ;
      RECT  6.910000  0.085000  7.170000 0.645000 ;
      RECT  7.770000  0.085000  8.030000 0.565000 ;
      RECT  8.630000  0.085000  8.890000 0.565000 ;
      RECT  9.490000  0.085000  9.735000 0.565000 ;
      RECT 10.350000  0.085000 10.595000 0.565000 ;
      RECT 11.205000  0.085000 11.455000 0.565000 ;
      RECT 12.065000  0.085000 12.315000 0.565000 ;
      RECT 12.925000  0.085000 13.185000 0.565000 ;
      RECT 13.785000  0.085000 14.085000 0.565000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.525000  0.765000  2.695000 0.935000 ;
      RECT  2.885000  0.765000  3.055000 0.935000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.210000  0.765000  5.380000 0.935000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
    LAYER met1 ;
      RECT 2.465000 0.735000 3.115000 0.780000 ;
      RECT 2.465000 0.780000 5.440000 0.920000 ;
      RECT 2.465000 0.920000 3.115000 0.965000 ;
      RECT 5.150000 0.735000 5.440000 0.780000 ;
      RECT 5.150000 0.920000 5.440000 0.965000 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrckapwr_16
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.070000 3.290000 1.540000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.402500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335000 0.290000 5.635000 0.980000 ;
        RECT 5.360000 0.980000 5.635000 2.370000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 6.440000 5.680000 ;
      LAYER pwell ;
        RECT 0.145000 4.595000 0.315000 5.120000 ;
        RECT 5.925000 4.595000 6.095000 5.120000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.500000 6.170000 3.640000 ;
        RECT 0.080000 3.455000 0.370000 3.500000 ;
        RECT 0.080000 3.640000 0.370000 3.685000 ;
        RECT 5.870000 3.455000 6.160000 3.500000 ;
        RECT 5.870000 3.640000 6.160000 3.685000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 4.135000 ;
        RECT  4.250000 1.305000 6.630000 4.135000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  PIN VPWRIN
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.380000 2.065000 2.390000 2.335000 ;
        RECT 2.060000 1.635000 2.390000 2.065000 ;
        RECT 2.060000 2.335000 2.390000 2.660000 ;
        RECT 2.060000 2.660000 2.810000 3.750000 ;
      LAYER mcon ;
        RECT 1.420000 2.115000 1.590000 2.285000 ;
        RECT 1.780000 2.115000 1.950000 2.285000 ;
        RECT 2.140000 2.115000 2.310000 2.285000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 6.170000 2.280000 ;
        RECT 1.360000 2.085000 2.370000 2.140000 ;
        RECT 1.360000 2.280000 2.370000 2.315000 ;
      LAYER nwell ;
        RECT 1.920000 1.305000 2.980000 4.135000 ;
    END
  END VPWRIN
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 1.890000 2.805000 ;
      RECT 0.000000  5.355000 6.440000 5.525000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  2.985000 0.375000 3.970000 ;
      RECT 0.085000  4.630000 0.375000 5.355000 ;
      RECT 2.020000  0.085000 2.350000 0.895000 ;
      RECT 2.560000  0.375000 2.800000 2.130000 ;
      RECT 2.560000  2.130000 3.390000 2.370000 ;
      RECT 2.645000  4.515000 2.905000 5.355000 ;
      RECT 3.060000  2.370000 3.390000 3.965000 ;
      RECT 3.075000  4.265000 4.265000 4.325000 ;
      RECT 3.075000  4.325000 3.405000 5.185000 ;
      RECT 3.115000  0.085000 3.445000 0.900000 ;
      RECT 3.145000  4.155000 4.195000 4.265000 ;
      RECT 3.575000  4.515000 3.765000 5.355000 ;
      RECT 3.615000  0.290000 3.805000 0.730000 ;
      RECT 3.615000  0.730000 4.665000 0.980000 ;
      RECT 3.680000  2.405000 4.190000 2.575000 ;
      RECT 3.680000  2.575000 3.850000 3.470000 ;
      RECT 3.680000  3.470000 4.720000 3.640000 ;
      RECT 3.935000  4.325000 4.265000 5.185000 ;
      RECT 3.975000  0.085000 4.305000 0.560000 ;
      RECT 4.020000  0.980000 4.190000 2.405000 ;
      RECT 4.020000  2.745000 4.640000 2.915000 ;
      RECT 4.020000  2.915000 4.190000 3.300000 ;
      RECT 4.020000  3.810000 4.190000 4.155000 ;
      RECT 4.390000  3.085000 4.720000 3.470000 ;
      RECT 4.410000  3.640000 4.720000 3.740000 ;
      RECT 4.445000  4.515000 4.955000 5.355000 ;
      RECT 4.470000  1.625000 4.640000 2.745000 ;
      RECT 4.475000  0.290000 4.665000 0.730000 ;
      RECT 4.835000  0.085000 5.165000 0.900000 ;
      RECT 4.890000  1.625000 5.120000 2.635000 ;
      RECT 4.890000  2.635000 6.440000 2.805000 ;
      RECT 4.890000  2.805000 5.120000 3.740000 ;
      RECT 5.135000  4.405000 5.765000 4.460000 ;
      RECT 5.135000  4.460000 5.695000 4.820000 ;
      RECT 5.135000  4.820000 5.485000 5.160000 ;
      RECT 5.360000  3.070000 5.550000 4.125000 ;
      RECT 5.360000  4.125000 6.085000 4.355000 ;
      RECT 5.360000  4.355000 5.765000 4.405000 ;
      RECT 5.865000  0.085000 6.155000 0.810000 ;
      RECT 5.865000  2.985000 6.155000 3.955000 ;
      RECT 5.865000  4.630000 6.155000 5.355000 ;
    LAYER mcon ;
      RECT 0.140000  3.485000 0.310000 3.655000 ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.145000  5.355000 0.315000 5.525000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.605000  5.355000 0.775000 5.525000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.065000  5.355000 1.235000 5.525000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.525000  5.355000 1.695000 5.525000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  5.355000 2.155000 5.525000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  5.355000 2.615000 5.525000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  5.355000 3.075000 5.525000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  5.355000 3.535000 5.525000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  5.355000 3.995000 5.525000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  5.355000 4.455000 5.525000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  5.355000 4.915000 5.525000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.205000  5.355000 5.375000 5.525000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.665000  5.355000 5.835000 5.525000 ;
      RECT 5.930000  3.485000 6.100000 3.655000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.125000  5.355000 6.295000 5.525000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 6.440000 0.240000 ;
    LAYER pwell ;
      RECT 0.145000 0.320000 0.315000 0.845000 ;
      RECT 5.925000 0.320000 6.095000 0.845000 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.070000 3.290000 1.540000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.610500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335000 0.255000 5.635000 0.980000 ;
        RECT 5.360000 0.980000 5.635000 2.370000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 6.440000 5.680000 ;
      LAYER pwell ;
        RECT 0.145000 4.595000 0.315000 5.120000 ;
        RECT 6.125000 4.595000 6.295000 5.120000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.500000 6.300000 3.640000 ;
        RECT 0.080000 3.455000 0.370000 3.500000 ;
        RECT 0.080000 3.640000 0.370000 3.685000 ;
        RECT 6.010000 3.455000 6.300000 3.500000 ;
        RECT 6.010000 3.640000 6.300000 3.685000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 4.135000 ;
        RECT  4.250000 1.305000 6.630000 4.135000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  PIN VPWRIN
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.380000 2.065000 2.390000 2.335000 ;
        RECT 2.060000 1.635000 2.390000 2.065000 ;
        RECT 2.060000 2.335000 2.390000 2.660000 ;
        RECT 2.060000 2.660000 2.810000 3.750000 ;
      LAYER mcon ;
        RECT 1.420000 2.115000 1.590000 2.285000 ;
        RECT 1.780000 2.115000 1.950000 2.285000 ;
        RECT 2.140000 2.115000 2.310000 2.285000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 6.370000 2.280000 ;
        RECT 1.360000 2.085000 2.370000 2.140000 ;
        RECT 1.360000 2.280000 2.370000 2.315000 ;
      LAYER nwell ;
        RECT 1.920000 1.305000 2.980000 4.135000 ;
    END
  END VPWRIN
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 1.890000 2.805000 ;
      RECT 0.000000  5.355000 6.440000 5.525000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  2.985000 0.375000 3.970000 ;
      RECT 0.085000  4.630000 0.375000 5.355000 ;
      RECT 2.020000  0.085000 2.350000 0.895000 ;
      RECT 2.560000  0.375000 2.800000 2.130000 ;
      RECT 2.560000  2.130000 3.390000 2.370000 ;
      RECT 2.645000  4.515000 2.905000 5.355000 ;
      RECT 3.060000  2.370000 3.390000 3.965000 ;
      RECT 3.075000  4.265000 4.265000 4.325000 ;
      RECT 3.075000  4.325000 3.405000 5.185000 ;
      RECT 3.115000  0.085000 3.445000 0.900000 ;
      RECT 3.145000  4.155000 4.195000 4.265000 ;
      RECT 3.575000  4.515000 3.765000 5.355000 ;
      RECT 3.615000  0.255000 3.805000 0.730000 ;
      RECT 3.615000  0.730000 4.665000 0.980000 ;
      RECT 3.680000  2.405000 4.190000 2.575000 ;
      RECT 3.680000  2.575000 3.850000 3.470000 ;
      RECT 3.680000  3.470000 4.720000 3.640000 ;
      RECT 3.935000  4.325000 4.265000 5.185000 ;
      RECT 3.975000  0.085000 4.305000 0.560000 ;
      RECT 4.020000  0.980000 4.190000 2.405000 ;
      RECT 4.020000  2.745000 4.640000 2.915000 ;
      RECT 4.020000  2.915000 4.190000 3.300000 ;
      RECT 4.020000  3.810000 4.190000 4.155000 ;
      RECT 4.390000  3.085000 4.720000 3.470000 ;
      RECT 4.410000  3.640000 4.720000 3.740000 ;
      RECT 4.445000  4.515000 4.955000 5.355000 ;
      RECT 4.470000  1.625000 4.640000 2.745000 ;
      RECT 4.475000  0.255000 4.665000 0.730000 ;
      RECT 4.835000  0.085000 5.165000 0.900000 ;
      RECT 4.890000  1.625000 5.120000 2.635000 ;
      RECT 4.890000  2.635000 6.440000 2.805000 ;
      RECT 4.890000  2.805000 5.120000 3.740000 ;
      RECT 5.135000  4.405000 5.765000 4.460000 ;
      RECT 5.135000  4.460000 5.695000 4.820000 ;
      RECT 5.135000  4.820000 5.485000 5.160000 ;
      RECT 5.360000  3.070000 5.550000 4.125000 ;
      RECT 5.360000  4.125000 6.085000 4.355000 ;
      RECT 5.360000  4.355000 5.765000 4.405000 ;
      RECT 5.825000  0.085000 6.155000 0.900000 ;
      RECT 5.905000  1.610000 6.075000 2.635000 ;
      RECT 6.065000  2.985000 6.355000 3.955000 ;
      RECT 6.065000  4.630000 6.355000 5.355000 ;
    LAYER mcon ;
      RECT 0.140000  3.485000 0.310000 3.655000 ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.145000  5.355000 0.315000 5.525000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.605000  5.355000 0.775000 5.525000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.065000  5.355000 1.235000 5.525000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.525000  5.355000 1.695000 5.525000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  5.355000 2.155000 5.525000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  5.355000 2.615000 5.525000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  5.355000 3.075000 5.525000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  5.355000 3.535000 5.525000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  5.355000 3.995000 5.525000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  5.355000 4.455000 5.525000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  5.355000 4.915000 5.525000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.205000  5.355000 5.375000 5.525000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.665000  5.355000 5.835000 5.525000 ;
      RECT 6.070000  3.485000 6.240000 3.655000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.125000  5.355000 6.295000 5.525000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 6.440000 0.240000 ;
    LAYER pwell ;
      RECT 0.145000 0.320000 0.315000 0.845000 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.070000 3.290000 1.540000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.072500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335000 0.255000 5.635000 0.980000 ;
        RECT 5.360000 0.980000 5.635000 1.085000 ;
        RECT 5.360000 1.085000 6.555000 1.410000 ;
        RECT 5.360000 1.410000 5.635000 2.370000 ;
        RECT 6.280000 1.410000 6.555000 2.370000 ;
        RECT 6.335000 0.255000 6.555000 1.085000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 7.360000 5.680000 ;
      LAYER pwell ;
        RECT 0.145000 4.595000 0.315000 5.120000 ;
        RECT 7.045000 4.595000 7.215000 5.120000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.500000 7.290000 3.640000 ;
        RECT 0.080000 3.455000 0.370000 3.500000 ;
        RECT 0.080000 3.640000 0.370000 3.685000 ;
        RECT 6.930000 3.455000 7.220000 3.500000 ;
        RECT 6.930000 3.640000 7.220000 3.685000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 4.135000 ;
        RECT  4.250000 1.305000 7.405000 4.135000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  PIN VPWRIN
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.380000 2.065000 2.390000 2.335000 ;
        RECT 2.060000 1.635000 2.390000 2.065000 ;
        RECT 2.060000 2.335000 2.390000 2.660000 ;
        RECT 2.060000 2.660000 2.810000 3.750000 ;
      LAYER mcon ;
        RECT 1.420000 2.115000 1.590000 2.285000 ;
        RECT 1.780000 2.115000 1.950000 2.285000 ;
        RECT 2.140000 2.115000 2.310000 2.285000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 7.290000 2.280000 ;
        RECT 1.360000 2.085000 2.370000 2.140000 ;
        RECT 1.360000 2.280000 2.370000 2.315000 ;
      LAYER nwell ;
        RECT 1.920000 1.305000 2.980000 4.135000 ;
    END
  END VPWRIN
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 1.890000 2.805000 ;
      RECT 0.000000  5.355000 7.360000 5.525000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  2.985000 0.375000 3.970000 ;
      RECT 0.085000  4.630000 0.375000 5.355000 ;
      RECT 2.020000  0.085000 2.350000 0.895000 ;
      RECT 2.560000  0.375000 2.800000 2.130000 ;
      RECT 2.560000  2.130000 3.390000 2.370000 ;
      RECT 2.645000  4.515000 2.905000 5.355000 ;
      RECT 3.060000  2.370000 3.390000 3.965000 ;
      RECT 3.075000  4.265000 4.265000 4.325000 ;
      RECT 3.075000  4.325000 3.405000 5.185000 ;
      RECT 3.115000  0.085000 3.445000 0.900000 ;
      RECT 3.145000  4.155000 4.195000 4.265000 ;
      RECT 3.575000  4.515000 3.765000 5.355000 ;
      RECT 3.615000  0.255000 3.805000 0.730000 ;
      RECT 3.615000  0.730000 4.665000 0.980000 ;
      RECT 3.680000  2.405000 4.190000 2.575000 ;
      RECT 3.680000  2.575000 3.850000 3.470000 ;
      RECT 3.680000  3.470000 4.720000 3.640000 ;
      RECT 3.935000  4.325000 4.265000 5.185000 ;
      RECT 3.975000  0.085000 4.305000 0.560000 ;
      RECT 4.020000  0.980000 4.190000 2.405000 ;
      RECT 4.020000  2.745000 4.640000 2.915000 ;
      RECT 4.020000  2.915000 4.190000 3.300000 ;
      RECT 4.020000  3.810000 4.190000 4.155000 ;
      RECT 4.390000  3.085000 4.720000 3.470000 ;
      RECT 4.410000  3.640000 4.720000 3.740000 ;
      RECT 4.445000  4.515000 4.955000 5.355000 ;
      RECT 4.470000  1.625000 4.640000 2.745000 ;
      RECT 4.475000  0.255000 4.665000 0.730000 ;
      RECT 4.835000  0.085000 5.165000 0.900000 ;
      RECT 4.890000  1.625000 5.120000 2.635000 ;
      RECT 4.890000  2.635000 7.360000 2.805000 ;
      RECT 4.890000  2.805000 5.120000 3.740000 ;
      RECT 5.135000  4.405000 5.765000 4.460000 ;
      RECT 5.135000  4.460000 5.695000 4.820000 ;
      RECT 5.135000  4.820000 5.485000 5.160000 ;
      RECT 5.360000  3.070000 5.550000 4.125000 ;
      RECT 5.360000  4.125000 6.085000 4.355000 ;
      RECT 5.360000  4.355000 5.765000 4.405000 ;
      RECT 5.825000  0.085000 6.155000 0.845000 ;
      RECT 5.905000  1.610000 6.075000 2.635000 ;
      RECT 6.755000  0.085000 7.005000 0.925000 ;
      RECT 6.755000  1.610000 6.935000 2.635000 ;
      RECT 6.985000  2.985000 7.275000 3.955000 ;
      RECT 6.985000  4.630000 7.275000 5.355000 ;
    LAYER mcon ;
      RECT 0.140000  3.485000 0.310000 3.655000 ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.145000  5.355000 0.315000 5.525000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.605000  5.355000 0.775000 5.525000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.065000  5.355000 1.235000 5.525000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.525000  5.355000 1.695000 5.525000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  5.355000 2.155000 5.525000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  5.355000 2.615000 5.525000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  5.355000 3.075000 5.525000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  5.355000 3.535000 5.525000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  5.355000 3.995000 5.525000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  5.355000 4.455000 5.525000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  5.355000 4.915000 5.525000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.205000  5.355000 5.375000 5.525000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.665000  5.355000 5.835000 5.525000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.125000  5.355000 6.295000 5.525000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.585000  5.355000 6.755000 5.525000 ;
      RECT 6.990000  3.485000 7.160000 3.655000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.045000  5.355000 7.215000 5.525000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 7.360000 0.240000 ;
    LAYER pwell ;
      RECT 0.145000 0.320000 0.315000 0.845000 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.070000 3.290000 1.540000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.072500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335000 0.255000 5.635000 0.980000 ;
        RECT 5.360000 0.980000 5.635000 1.085000 ;
        RECT 5.360000 1.085000 6.555000 1.410000 ;
        RECT 5.360000 1.410000 5.635000 2.370000 ;
        RECT 6.280000 1.410000 6.555000 2.370000 ;
        RECT 6.335000 0.255000 6.555000 1.085000 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.380000 2.065000 2.390000 2.335000 ;
        RECT 2.060000 1.635000 2.390000 2.065000 ;
        RECT 2.060000 2.335000 2.390000 2.660000 ;
        RECT 2.060000 2.660000 2.810000 3.750000 ;
      LAYER mcon ;
        RECT 1.420000 2.115000 1.590000 2.285000 ;
        RECT 1.780000 2.115000 1.950000 2.285000 ;
        RECT 2.140000 2.115000 2.310000 2.285000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 7.290000 2.280000 ;
        RECT 1.360000 2.085000 2.370000 2.140000 ;
        RECT 1.360000 2.280000 2.370000 2.315000 ;
      LAYER nwell ;
        RECT 1.920000 1.305000 2.980000 4.135000 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 7.360000 5.680000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.075000 5.245000 0.200000 5.395000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 4.250000 1.305000 7.405000 4.135000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 1.890000 2.805000 ;
      RECT 0.000000  5.355000 7.360000 5.525000 ;
      RECT 2.020000  0.085000 2.350000 0.895000 ;
      RECT 2.560000  0.375000 2.800000 2.130000 ;
      RECT 2.560000  2.130000 3.390000 2.370000 ;
      RECT 2.645000  4.515000 2.905000 5.355000 ;
      RECT 3.060000  2.370000 3.390000 3.965000 ;
      RECT 3.075000  4.265000 4.265000 4.325000 ;
      RECT 3.075000  4.325000 3.405000 5.185000 ;
      RECT 3.115000  0.085000 3.445000 0.900000 ;
      RECT 3.145000  4.155000 4.195000 4.265000 ;
      RECT 3.575000  4.515000 3.765000 5.355000 ;
      RECT 3.615000  0.255000 3.805000 0.730000 ;
      RECT 3.615000  0.730000 4.665000 0.980000 ;
      RECT 3.680000  2.405000 4.190000 2.575000 ;
      RECT 3.680000  2.575000 3.850000 3.470000 ;
      RECT 3.680000  3.470000 4.720000 3.640000 ;
      RECT 3.935000  4.325000 4.265000 5.185000 ;
      RECT 3.975000  0.085000 4.305000 0.560000 ;
      RECT 4.020000  0.980000 4.190000 2.405000 ;
      RECT 4.020000  2.745000 4.640000 2.915000 ;
      RECT 4.020000  2.915000 4.190000 3.300000 ;
      RECT 4.020000  3.810000 4.190000 4.155000 ;
      RECT 4.390000  3.085000 4.720000 3.470000 ;
      RECT 4.410000  3.640000 4.720000 3.740000 ;
      RECT 4.445000  4.515000 4.955000 5.355000 ;
      RECT 4.470000  1.625000 4.640000 2.745000 ;
      RECT 4.475000  0.255000 4.665000 0.730000 ;
      RECT 4.835000  0.085000 5.165000 0.900000 ;
      RECT 4.890000  1.625000 5.120000 2.635000 ;
      RECT 4.890000  2.635000 7.360000 2.805000 ;
      RECT 4.890000  2.805000 5.120000 3.740000 ;
      RECT 5.135000  4.405000 5.765000 4.460000 ;
      RECT 5.135000  4.460000 5.695000 4.820000 ;
      RECT 5.135000  4.820000 5.485000 5.160000 ;
      RECT 5.360000  3.070000 5.550000 4.125000 ;
      RECT 5.360000  4.125000 6.085000 4.355000 ;
      RECT 5.360000  4.355000 5.765000 4.405000 ;
      RECT 5.825000  0.085000 6.155000 0.845000 ;
      RECT 5.905000  1.610000 6.075000 2.635000 ;
      RECT 6.755000  0.085000 7.005000 0.925000 ;
      RECT 6.755000  1.610000 6.935000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.145000  5.355000 0.315000 5.525000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.605000  5.355000 0.775000 5.525000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.065000  5.355000 1.235000 5.525000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.525000  5.355000 1.695000 5.525000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  5.355000 2.155000 5.525000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  5.355000 2.615000 5.525000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  5.355000 3.075000 5.525000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  5.355000 3.535000 5.525000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  5.355000 3.995000 5.525000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  5.355000 4.455000 5.525000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  5.355000 4.915000 5.525000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.205000  5.355000 5.375000 5.525000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.665000  5.355000 5.835000 5.525000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.125000  5.355000 6.295000 5.525000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.585000  5.355000 6.755000 5.525000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.045000  5.355000 7.215000 5.525000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 7.360000 0.240000 ;
    LAYER nwell ;
      RECT -0.190000 1.305000 0.650000 4.135000 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.070000 3.290000 1.540000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.402500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335000 0.290000 5.635000 0.980000 ;
        RECT 5.360000 0.980000 5.635000 2.370000 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.380000 2.065000 2.390000 2.335000 ;
        RECT 2.060000 1.635000 2.390000 2.065000 ;
        RECT 2.060000 2.335000 2.390000 2.660000 ;
        RECT 2.060000 2.660000 2.810000 3.750000 ;
      LAYER mcon ;
        RECT 1.420000 2.115000 1.590000 2.285000 ;
        RECT 1.780000 2.115000 1.950000 2.285000 ;
        RECT 2.140000 2.115000 2.310000 2.285000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 6.170000 2.280000 ;
        RECT 1.360000 2.085000 2.370000 2.140000 ;
        RECT 1.360000 2.280000 2.370000 2.315000 ;
      LAYER nwell ;
        RECT 1.920000 1.305000 2.980000 4.135000 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 6.440000 5.680000 ;
      LAYER pwell ;
        RECT 0.145000 4.595000 0.315000 5.120000 ;
        RECT 5.925000 4.595000 6.095000 5.120000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.500000 6.170000 3.640000 ;
        RECT 0.080000 3.455000 0.370000 3.500000 ;
        RECT 0.080000 3.640000 0.370000 3.685000 ;
        RECT 5.870000 3.455000 6.160000 3.500000 ;
        RECT 5.870000 3.640000 6.160000 3.685000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 4.135000 ;
        RECT  4.250000 1.305000 6.630000 4.135000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 1.890000 2.805000 ;
      RECT 0.000000  5.355000 6.440000 5.525000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  2.985000 0.375000 3.970000 ;
      RECT 0.085000  4.630000 0.375000 5.355000 ;
      RECT 2.020000  0.085000 2.350000 0.895000 ;
      RECT 2.560000  0.375000 2.800000 2.130000 ;
      RECT 2.560000  2.130000 3.390000 2.370000 ;
      RECT 2.645000  4.515000 2.905000 5.355000 ;
      RECT 3.060000  2.370000 3.390000 3.965000 ;
      RECT 3.075000  4.265000 4.265000 4.325000 ;
      RECT 3.075000  4.325000 3.405000 5.185000 ;
      RECT 3.115000  0.085000 3.445000 0.900000 ;
      RECT 3.145000  4.155000 4.195000 4.265000 ;
      RECT 3.575000  4.515000 3.765000 5.355000 ;
      RECT 3.615000  0.290000 3.805000 0.730000 ;
      RECT 3.615000  0.730000 4.665000 0.980000 ;
      RECT 3.680000  2.405000 4.190000 2.575000 ;
      RECT 3.680000  2.575000 3.850000 3.470000 ;
      RECT 3.680000  3.470000 4.720000 3.640000 ;
      RECT 3.935000  4.325000 4.265000 5.185000 ;
      RECT 3.975000  0.085000 4.305000 0.560000 ;
      RECT 4.020000  0.980000 4.190000 2.405000 ;
      RECT 4.020000  2.745000 4.640000 2.915000 ;
      RECT 4.020000  2.915000 4.190000 3.300000 ;
      RECT 4.020000  3.810000 4.190000 4.155000 ;
      RECT 4.390000  3.085000 4.720000 3.470000 ;
      RECT 4.410000  3.640000 4.720000 3.740000 ;
      RECT 4.445000  4.515000 4.955000 5.355000 ;
      RECT 4.470000  1.625000 4.640000 2.745000 ;
      RECT 4.475000  0.290000 4.665000 0.730000 ;
      RECT 4.835000  0.085000 5.165000 0.900000 ;
      RECT 4.890000  1.625000 5.120000 2.635000 ;
      RECT 4.890000  2.635000 6.440000 2.805000 ;
      RECT 4.890000  2.805000 5.120000 3.740000 ;
      RECT 5.135000  4.405000 5.765000 4.460000 ;
      RECT 5.135000  4.460000 5.695000 4.820000 ;
      RECT 5.135000  4.820000 5.485000 5.160000 ;
      RECT 5.360000  3.070000 5.550000 4.125000 ;
      RECT 5.360000  4.125000 6.085000 4.355000 ;
      RECT 5.360000  4.355000 5.765000 4.405000 ;
      RECT 5.865000  0.085000 6.155000 0.810000 ;
      RECT 5.865000  2.985000 6.155000 3.955000 ;
      RECT 5.865000  4.630000 6.155000 5.355000 ;
    LAYER mcon ;
      RECT 0.140000  3.485000 0.310000 3.655000 ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.145000  5.355000 0.315000 5.525000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.605000  5.355000 0.775000 5.525000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.065000  5.355000 1.235000 5.525000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.525000  5.355000 1.695000 5.525000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  5.355000 2.155000 5.525000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  5.355000 2.615000 5.525000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  5.355000 3.075000 5.525000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  5.355000 3.535000 5.525000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  5.355000 3.995000 5.525000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  5.355000 4.455000 5.525000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  5.355000 4.915000 5.525000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.205000  5.355000 5.375000 5.525000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.665000  5.355000 5.835000 5.525000 ;
      RECT 5.930000  3.485000 6.100000 3.655000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.125000  5.355000 6.295000 5.525000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 6.440000 0.240000 ;
    LAYER pwell ;
      RECT 0.145000 0.320000 0.315000 0.845000 ;
      RECT 5.925000 0.320000 6.095000 0.845000 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.070000 3.290000 1.540000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.610500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335000 0.255000 5.635000 0.980000 ;
        RECT 5.360000 0.980000 5.635000 2.370000 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.380000 2.065000 2.390000 2.335000 ;
        RECT 2.060000 1.635000 2.390000 2.065000 ;
        RECT 2.060000 2.335000 2.390000 2.660000 ;
        RECT 2.060000 2.660000 2.810000 3.750000 ;
      LAYER mcon ;
        RECT 1.420000 2.115000 1.590000 2.285000 ;
        RECT 1.780000 2.115000 1.950000 2.285000 ;
        RECT 2.140000 2.115000 2.310000 2.285000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 6.370000 2.280000 ;
        RECT 1.360000 2.085000 2.370000 2.140000 ;
        RECT 1.360000 2.280000 2.370000 2.315000 ;
      LAYER nwell ;
        RECT 1.920000 1.305000 2.980000 4.135000 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 6.440000 5.680000 ;
      LAYER pwell ;
        RECT 0.145000 4.595000 0.315000 5.120000 ;
        RECT 6.125000 4.595000 6.295000 5.120000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.500000 6.300000 3.640000 ;
        RECT 0.080000 3.455000 0.370000 3.500000 ;
        RECT 0.080000 3.640000 0.370000 3.685000 ;
        RECT 6.010000 3.455000 6.300000 3.500000 ;
        RECT 6.010000 3.640000 6.300000 3.685000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 4.135000 ;
        RECT  4.250000 1.305000 6.630000 4.135000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 1.890000 2.805000 ;
      RECT 0.000000  5.355000 6.440000 5.525000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  2.985000 0.375000 3.970000 ;
      RECT 0.085000  4.630000 0.375000 5.355000 ;
      RECT 2.020000  0.085000 2.350000 0.895000 ;
      RECT 2.560000  0.375000 2.800000 2.130000 ;
      RECT 2.560000  2.130000 3.390000 2.370000 ;
      RECT 2.645000  4.515000 2.905000 5.355000 ;
      RECT 3.060000  2.370000 3.390000 3.965000 ;
      RECT 3.075000  4.265000 4.265000 4.325000 ;
      RECT 3.075000  4.325000 3.405000 5.185000 ;
      RECT 3.115000  0.085000 3.445000 0.900000 ;
      RECT 3.145000  4.155000 4.195000 4.265000 ;
      RECT 3.575000  4.515000 3.765000 5.355000 ;
      RECT 3.615000  0.255000 3.805000 0.730000 ;
      RECT 3.615000  0.730000 4.665000 0.980000 ;
      RECT 3.680000  2.405000 4.190000 2.575000 ;
      RECT 3.680000  2.575000 3.850000 3.470000 ;
      RECT 3.680000  3.470000 4.720000 3.640000 ;
      RECT 3.935000  4.325000 4.265000 5.185000 ;
      RECT 3.975000  0.085000 4.305000 0.560000 ;
      RECT 4.020000  0.980000 4.190000 2.405000 ;
      RECT 4.020000  2.745000 4.640000 2.915000 ;
      RECT 4.020000  2.915000 4.190000 3.300000 ;
      RECT 4.020000  3.810000 4.190000 4.155000 ;
      RECT 4.390000  3.085000 4.720000 3.470000 ;
      RECT 4.410000  3.640000 4.720000 3.740000 ;
      RECT 4.445000  4.515000 4.955000 5.355000 ;
      RECT 4.470000  1.625000 4.640000 2.745000 ;
      RECT 4.475000  0.255000 4.665000 0.730000 ;
      RECT 4.835000  0.085000 5.165000 0.900000 ;
      RECT 4.890000  1.625000 5.120000 2.635000 ;
      RECT 4.890000  2.635000 6.440000 2.805000 ;
      RECT 4.890000  2.805000 5.120000 3.740000 ;
      RECT 5.135000  4.405000 5.765000 4.460000 ;
      RECT 5.135000  4.460000 5.695000 4.820000 ;
      RECT 5.135000  4.820000 5.485000 5.160000 ;
      RECT 5.360000  3.070000 5.550000 4.125000 ;
      RECT 5.360000  4.125000 6.085000 4.355000 ;
      RECT 5.360000  4.355000 5.765000 4.405000 ;
      RECT 5.825000  0.085000 6.155000 0.900000 ;
      RECT 5.905000  1.610000 6.075000 2.635000 ;
      RECT 6.065000  2.985000 6.355000 3.955000 ;
      RECT 6.065000  4.630000 6.355000 5.355000 ;
    LAYER mcon ;
      RECT 0.140000  3.485000 0.310000 3.655000 ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.145000  5.355000 0.315000 5.525000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.605000  5.355000 0.775000 5.525000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.065000  5.355000 1.235000 5.525000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.525000  5.355000 1.695000 5.525000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  5.355000 2.155000 5.525000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  5.355000 2.615000 5.525000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  5.355000 3.075000 5.525000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  5.355000 3.535000 5.525000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  5.355000 3.995000 5.525000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  5.355000 4.455000 5.525000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  5.355000 4.915000 5.525000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.205000  5.355000 5.375000 5.525000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.665000  5.355000 5.835000 5.525000 ;
      RECT 6.070000  3.485000 6.240000 3.655000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.125000  5.355000 6.295000 5.525000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 6.440000 0.240000 ;
    LAYER pwell ;
      RECT 0.145000 0.320000 0.315000 0.845000 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.070000 3.290000 1.540000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.072500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335000 0.255000 5.635000 0.980000 ;
        RECT 5.360000 0.980000 5.635000 1.085000 ;
        RECT 5.360000 1.085000 6.555000 1.410000 ;
        RECT 5.360000 1.410000 5.635000 2.370000 ;
        RECT 6.280000 1.410000 6.555000 2.370000 ;
        RECT 6.335000 0.255000 6.555000 1.085000 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.380000 2.065000 2.390000 2.335000 ;
        RECT 2.060000 1.635000 2.390000 2.065000 ;
        RECT 2.060000 2.335000 2.390000 2.660000 ;
        RECT 2.060000 2.660000 2.810000 3.750000 ;
      LAYER mcon ;
        RECT 1.420000 2.115000 1.590000 2.285000 ;
        RECT 1.780000 2.115000 1.950000 2.285000 ;
        RECT 2.140000 2.115000 2.310000 2.285000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 7.290000 2.280000 ;
        RECT 1.360000 2.085000 2.370000 2.140000 ;
        RECT 1.360000 2.280000 2.370000 2.315000 ;
      LAYER nwell ;
        RECT 1.920000 1.305000 2.980000 4.135000 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 7.360000 5.680000 ;
      LAYER pwell ;
        RECT 0.145000 4.595000 0.315000 5.120000 ;
        RECT 7.045000 4.595000 7.215000 5.120000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.500000 7.290000 3.640000 ;
        RECT 0.080000 3.455000 0.370000 3.500000 ;
        RECT 0.080000 3.640000 0.370000 3.685000 ;
        RECT 6.930000 3.455000 7.220000 3.500000 ;
        RECT 6.930000 3.640000 7.220000 3.685000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 4.135000 ;
        RECT  4.250000 1.305000 7.405000 4.135000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 1.890000 2.805000 ;
      RECT 0.000000  5.355000 7.360000 5.525000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  2.985000 0.375000 3.970000 ;
      RECT 0.085000  4.630000 0.375000 5.355000 ;
      RECT 2.020000  0.085000 2.350000 0.895000 ;
      RECT 2.560000  0.375000 2.800000 2.130000 ;
      RECT 2.560000  2.130000 3.390000 2.370000 ;
      RECT 2.645000  4.515000 2.905000 5.355000 ;
      RECT 3.060000  2.370000 3.390000 3.965000 ;
      RECT 3.075000  4.265000 4.265000 4.325000 ;
      RECT 3.075000  4.325000 3.405000 5.185000 ;
      RECT 3.115000  0.085000 3.445000 0.900000 ;
      RECT 3.145000  4.155000 4.195000 4.265000 ;
      RECT 3.575000  4.515000 3.765000 5.355000 ;
      RECT 3.615000  0.255000 3.805000 0.730000 ;
      RECT 3.615000  0.730000 4.665000 0.980000 ;
      RECT 3.680000  2.405000 4.190000 2.575000 ;
      RECT 3.680000  2.575000 3.850000 3.470000 ;
      RECT 3.680000  3.470000 4.720000 3.640000 ;
      RECT 3.935000  4.325000 4.265000 5.185000 ;
      RECT 3.975000  0.085000 4.305000 0.560000 ;
      RECT 4.020000  0.980000 4.190000 2.405000 ;
      RECT 4.020000  2.745000 4.640000 2.915000 ;
      RECT 4.020000  2.915000 4.190000 3.300000 ;
      RECT 4.020000  3.810000 4.190000 4.155000 ;
      RECT 4.390000  3.085000 4.720000 3.470000 ;
      RECT 4.410000  3.640000 4.720000 3.740000 ;
      RECT 4.445000  4.515000 4.955000 5.355000 ;
      RECT 4.470000  1.625000 4.640000 2.745000 ;
      RECT 4.475000  0.255000 4.665000 0.730000 ;
      RECT 4.835000  0.085000 5.165000 0.900000 ;
      RECT 4.890000  1.625000 5.120000 2.635000 ;
      RECT 4.890000  2.635000 7.360000 2.805000 ;
      RECT 4.890000  2.805000 5.120000 3.740000 ;
      RECT 5.135000  4.405000 5.765000 4.460000 ;
      RECT 5.135000  4.460000 5.695000 4.820000 ;
      RECT 5.135000  4.820000 5.485000 5.160000 ;
      RECT 5.360000  3.070000 5.550000 4.125000 ;
      RECT 5.360000  4.125000 6.085000 4.355000 ;
      RECT 5.360000  4.355000 5.765000 4.405000 ;
      RECT 5.825000  0.085000 6.155000 0.845000 ;
      RECT 5.905000  1.610000 6.075000 2.635000 ;
      RECT 6.755000  0.085000 7.005000 0.925000 ;
      RECT 6.755000  1.610000 6.935000 2.635000 ;
      RECT 6.985000  2.985000 7.275000 3.955000 ;
      RECT 6.985000  4.630000 7.275000 5.355000 ;
    LAYER mcon ;
      RECT 0.140000  3.485000 0.310000 3.655000 ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.145000  5.355000 0.315000 5.525000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.605000  5.355000 0.775000 5.525000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.065000  5.355000 1.235000 5.525000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.525000  5.355000 1.695000 5.525000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  5.355000 2.155000 5.525000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  5.355000 2.615000 5.525000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  5.355000 3.075000 5.525000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  5.355000 3.535000 5.525000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  5.355000 3.995000 5.525000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  5.355000 4.455000 5.525000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  5.355000 4.915000 5.525000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.205000  5.355000 5.375000 5.525000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.665000  5.355000 5.835000 5.525000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.125000  5.355000 6.295000 5.525000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.585000  5.355000 6.755000 5.525000 ;
      RECT 6.990000  3.485000 7.160000 3.655000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.045000  5.355000 7.215000 5.525000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 7.360000 0.240000 ;
    LAYER pwell ;
      RECT 0.145000 0.320000 0.315000 0.845000 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4
MACRO sky130_fd_sc_hd__macro_sparecell
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__macro_sparecell ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.34000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN LO
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.215000 1.075000 4.965000 1.325000 ;
      LAYER mcon ;
        RECT 4.775000 1.105000 4.945000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.135000 1.075000 5.895000 1.325000 ;
      LAYER mcon ;
        RECT 5.705000 1.105000 5.875000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.755000 0.915000 7.275000 2.465000 ;
      LAYER mcon ;
        RECT 6.765000 1.105000 6.935000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.445000 1.075000 8.205000 1.325000 ;
      LAYER mcon ;
        RECT 7.625000 1.105000 7.795000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.375000 1.075000 9.125000 1.325000 ;
      LAYER mcon ;
        RECT 8.485000 1.105000 8.655000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.715000 1.075000 5.005000 1.120000 ;
        RECT 4.715000 1.120000 8.715000 1.260000 ;
        RECT 4.715000 1.260000 5.005000 1.305000 ;
        RECT 5.645000 1.075000 5.935000 1.120000 ;
        RECT 5.645000 1.260000 5.935000 1.305000 ;
        RECT 6.705000 1.075000 6.995000 1.120000 ;
        RECT 6.705000 1.260000 6.995000 1.305000 ;
        RECT 7.565000 1.075000 7.855000 1.120000 ;
        RECT 7.565000 1.260000 7.855000 1.305000 ;
        RECT 8.425000 1.075000 8.715000 1.120000 ;
        RECT 8.425000 1.260000 8.715000 1.305000 ;
    END
  END LO
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 13.340000 0.085000 ;
        RECT  0.145000  0.085000  0.355000 0.905000 ;
        RECT  1.025000  0.085000  1.255000 0.905000 ;
        RECT  1.515000  0.085000  1.805000 0.555000 ;
        RECT  2.475000  0.085000  2.645000 0.555000 ;
        RECT  3.315000  0.085000  3.590000 0.905000 ;
        RECT  5.215000  0.085000  5.385000 0.545000 ;
        RECT  6.755000  0.085000  7.095000 0.745000 ;
        RECT  7.955000  0.085000  8.125000 0.545000 ;
        RECT  9.750000  0.085000 10.025000 0.905000 ;
        RECT 10.695000  0.085000 10.865000 0.555000 ;
        RECT 11.535000  0.085000 11.825000 0.555000 ;
        RECT 12.085000  0.085000 12.315000 0.905000 ;
        RECT 12.985000  0.085000 13.195000 0.905000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
        RECT 10.725000 -0.085000 10.895000 0.085000 ;
        RECT 11.185000 -0.085000 11.355000 0.085000 ;
        RECT 11.645000 -0.085000 11.815000 0.085000 ;
        RECT 12.105000 -0.085000 12.275000 0.085000 ;
        RECT 12.565000 -0.085000 12.735000 0.085000 ;
        RECT 13.025000 -0.085000 13.195000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.340000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 13.530000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 13.340000 2.805000 ;
        RECT  0.145000 1.495000  0.355000 2.635000 ;
        RECT  1.025000 1.495000  1.255000 2.635000 ;
        RECT  2.815000 1.835000  3.145000 2.635000 ;
        RECT  3.870000 1.835000  4.125000 2.635000 ;
        RECT  4.795000 1.835000  4.965000 2.635000 ;
        RECT  5.635000 1.495000  5.895000 2.635000 ;
        RECT  6.255000 1.910000  6.585000 2.635000 ;
        RECT  7.445000 1.495000  7.705000 2.635000 ;
        RECT  8.375000 1.835000  8.545000 2.635000 ;
        RECT  9.215000 1.835000  9.470000 2.635000 ;
        RECT 10.195000 1.835000 10.525000 2.635000 ;
        RECT 12.085000 1.495000 12.315000 2.635000 ;
        RECT 12.985000 1.495000 13.195000 2.635000 ;
      LAYER mcon ;
        RECT  0.145000 2.635000  0.315000 2.805000 ;
        RECT  0.605000 2.635000  0.775000 2.805000 ;
        RECT  1.065000 2.635000  1.235000 2.805000 ;
        RECT  1.525000 2.635000  1.695000 2.805000 ;
        RECT  1.985000 2.635000  2.155000 2.805000 ;
        RECT  2.445000 2.635000  2.615000 2.805000 ;
        RECT  2.905000 2.635000  3.075000 2.805000 ;
        RECT  3.365000 2.635000  3.535000 2.805000 ;
        RECT  3.825000 2.635000  3.995000 2.805000 ;
        RECT  4.285000 2.635000  4.455000 2.805000 ;
        RECT  4.745000 2.635000  4.915000 2.805000 ;
        RECT  5.205000 2.635000  5.375000 2.805000 ;
        RECT  5.665000 2.635000  5.835000 2.805000 ;
        RECT  6.125000 2.635000  6.295000 2.805000 ;
        RECT  6.585000 2.635000  6.755000 2.805000 ;
        RECT  7.045000 2.635000  7.215000 2.805000 ;
        RECT  7.505000 2.635000  7.675000 2.805000 ;
        RECT  7.965000 2.635000  8.135000 2.805000 ;
        RECT  8.425000 2.635000  8.595000 2.805000 ;
        RECT  8.885000 2.635000  9.055000 2.805000 ;
        RECT  9.345000 2.635000  9.515000 2.805000 ;
        RECT  9.805000 2.635000  9.975000 2.805000 ;
        RECT 10.265000 2.635000 10.435000 2.805000 ;
        RECT 10.725000 2.635000 10.895000 2.805000 ;
        RECT 11.185000 2.635000 11.355000 2.805000 ;
        RECT 11.645000 2.635000 11.815000 2.805000 ;
        RECT 12.105000 2.635000 12.275000 2.805000 ;
        RECT 12.565000 2.635000 12.735000 2.805000 ;
        RECT 13.025000 2.635000 13.195000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.340000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.525000 0.255000  0.855000 0.885000 ;
      RECT  0.525000 0.885000  0.775000 1.485000 ;
      RECT  0.525000 1.485000  0.855000 2.465000 ;
      RECT  0.945000 1.075000  1.275000 1.325000 ;
      RECT  1.505000 1.835000  1.805000 2.295000 ;
      RECT  1.505000 2.295000  2.645000 2.465000 ;
      RECT  1.545000 0.735000  3.145000 0.905000 ;
      RECT  1.545000 0.905000  1.760000 1.445000 ;
      RECT  1.545000 1.445000  2.305000 1.665000 ;
      RECT  1.930000 1.075000  2.700000 1.275000 ;
      RECT  1.975000 0.255000  2.305000 0.725000 ;
      RECT  1.975000 0.725000  3.145000 0.735000 ;
      RECT  1.975000 1.665000  2.305000 2.125000 ;
      RECT  2.475000 1.455000  3.590000 1.665000 ;
      RECT  2.475000 1.665000  2.645000 2.295000 ;
      RECT  2.815000 0.255000  3.145000 0.725000 ;
      RECT  2.870000 1.075000  3.590000 1.275000 ;
      RECT  3.315000 1.665000  3.590000 2.465000 ;
      RECT  3.765000 0.655000  4.625000 0.905000 ;
      RECT  3.765000 0.905000  4.045000 1.495000 ;
      RECT  3.765000 1.495000  5.465000 1.665000 ;
      RECT  3.875000 0.255000  5.045000 0.465000 ;
      RECT  3.875000 0.465000  4.205000 0.485000 ;
      RECT  4.295000 1.665000  4.625000 2.465000 ;
      RECT  4.795000 0.465000  5.045000 0.715000 ;
      RECT  4.795000 0.715000  5.895000 0.885000 ;
      RECT  5.135000 1.665000  5.465000 2.465000 ;
      RECT  5.555000 0.255000  5.895000 0.715000 ;
      RECT  6.065000 0.255000  6.585000 1.740000 ;
      RECT  7.445000 0.255000  7.785000 0.715000 ;
      RECT  7.445000 0.715000  8.545000 0.885000 ;
      RECT  7.875000 1.495000  9.575000 1.665000 ;
      RECT  7.875000 1.665000  8.205000 2.465000 ;
      RECT  8.295000 0.255000  9.465000 0.465000 ;
      RECT  8.295000 0.465000  8.545000 0.715000 ;
      RECT  8.715000 0.655000  9.575000 0.905000 ;
      RECT  8.715000 1.665000  9.045000 2.465000 ;
      RECT  9.135000 0.465000  9.465000 0.485000 ;
      RECT  9.295000 0.905000  9.575000 1.495000 ;
      RECT  9.750000 1.075000 10.470000 1.275000 ;
      RECT  9.750000 1.455000 10.865000 1.665000 ;
      RECT  9.750000 1.665000 10.025000 2.465000 ;
      RECT 10.195000 0.255000 10.525000 0.725000 ;
      RECT 10.195000 0.725000 11.365000 0.735000 ;
      RECT 10.195000 0.735000 11.795000 0.905000 ;
      RECT 10.640000 1.075000 11.410000 1.275000 ;
      RECT 10.695000 1.665000 10.865000 2.295000 ;
      RECT 10.695000 2.295000 11.835000 2.465000 ;
      RECT 11.035000 0.255000 11.365000 0.725000 ;
      RECT 11.035000 1.445000 11.795000 1.665000 ;
      RECT 11.035000 1.665000 11.365000 2.125000 ;
      RECT 11.535000 1.835000 11.835000 2.295000 ;
      RECT 11.580000 0.905000 11.795000 1.445000 ;
      RECT 12.065000 1.075000 12.395000 1.325000 ;
      RECT 12.485000 0.255000 12.815000 0.885000 ;
      RECT 12.485000 1.485000 12.815000 2.465000 ;
      RECT 12.565000 0.885000 12.815000 1.485000 ;
    LAYER mcon ;
      RECT  0.565000 1.105000  0.735000 1.275000 ;
      RECT  1.085000 1.105000  1.255000 1.275000 ;
      RECT  1.570000 1.105000  1.740000 1.275000 ;
      RECT  2.100000 1.105000  2.270000 1.275000 ;
      RECT  2.960000 1.105000  3.130000 1.275000 ;
      RECT  3.820000 1.105000  3.990000 1.275000 ;
      RECT  9.345000 1.105000  9.515000 1.275000 ;
      RECT 10.205000 1.105000 10.375000 1.275000 ;
      RECT 11.065000 1.105000 11.235000 1.275000 ;
      RECT 11.605000 1.105000 11.775000 1.275000 ;
      RECT 12.090000 1.105000 12.260000 1.275000 ;
      RECT 12.605000 1.105000 12.775000 1.275000 ;
    LAYER met1 ;
      RECT  0.505000 1.075000  0.875000 1.305000 ;
      RECT  1.025000 1.075000  1.315000 1.120000 ;
      RECT  1.025000 1.120000  1.800000 1.260000 ;
      RECT  1.025000 1.260000  1.315000 1.305000 ;
      RECT  1.510000 1.075000  1.800000 1.120000 ;
      RECT  1.510000 1.260000  1.800000 1.305000 ;
      RECT  2.040000 1.075000  2.330000 1.120000 ;
      RECT  2.040000 1.120000  4.050000 1.260000 ;
      RECT  2.040000 1.260000  2.330000 1.305000 ;
      RECT  2.900000 1.075000  3.190000 1.120000 ;
      RECT  2.900000 1.260000  3.190000 1.305000 ;
      RECT  3.760000 1.075000  4.050000 1.120000 ;
      RECT  3.760000 1.260000  4.050000 1.305000 ;
      RECT  9.285000 1.075000  9.575000 1.120000 ;
      RECT  9.285000 1.120000 11.295000 1.260000 ;
      RECT  9.285000 1.260000  9.575000 1.305000 ;
      RECT 10.145000 1.075000 10.435000 1.120000 ;
      RECT 10.145000 1.260000 10.435000 1.305000 ;
      RECT 11.005000 1.075000 11.295000 1.120000 ;
      RECT 11.005000 1.260000 11.295000 1.305000 ;
      RECT 11.545000 1.075000 11.835000 1.120000 ;
      RECT 11.545000 1.120000 12.320000 1.260000 ;
      RECT 11.545000 1.260000 11.835000 1.305000 ;
      RECT 12.030000 1.075000 12.320000 1.120000 ;
      RECT 12.030000 1.260000 12.320000 1.305000 ;
      RECT 12.470000 1.075000 12.835000 1.305000 ;
    LAYER pwell ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  3.360000 -0.085000  3.530000 0.085000 ;
      RECT  5.660000 -0.085000  5.830000 0.085000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  7.510000 -0.085000  7.680000 0.085000 ;
      RECT  9.810000 -0.085000  9.980000 0.085000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
  END
END sky130_fd_sc_hd__macro_sparecell
MACRO sky130_fd_sc_hd__maj3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__maj3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 0.995000 1.125000 1.325000 ;
        RECT 0.610000 1.325000 0.780000 2.460000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 0.995000 1.905000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415000 0.765000 2.755000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.602250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.255000 0.255000 3.595000 0.825000 ;
        RECT 3.255000 2.160000 3.595000 2.465000 ;
        RECT 3.265000 1.495000 3.595000 2.160000 ;
        RECT 3.370000 0.825000 3.595000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.135000  0.255000 0.395000 0.655000 ;
      RECT 0.135000  0.655000 2.245000 0.825000 ;
      RECT 0.135000  0.825000 0.395000 2.125000 ;
      RECT 0.875000  0.085000 1.205000 0.485000 ;
      RECT 0.955000  1.715000 1.205000 2.635000 ;
      RECT 1.655000  0.255000 1.985000 0.640000 ;
      RECT 1.655000  0.640000 2.245000 0.655000 ;
      RECT 1.655000  1.815000 2.245000 2.080000 ;
      RECT 2.075000  0.825000 2.245000 1.495000 ;
      RECT 2.075000  1.495000 3.095000 1.665000 ;
      RECT 2.075000  1.665000 2.245000 1.815000 ;
      RECT 2.545000  0.085000 2.880000 0.470000 ;
      RECT 2.555000  1.845000 2.885000 2.635000 ;
      RECT 2.925000  0.995000 3.200000 1.325000 ;
      RECT 2.925000  1.325000 3.095000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__maj3_1
MACRO sky130_fd_sc_hd__maj3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__maj3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 0.995000 1.695000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.865000 0.995000 2.155000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.495000 ;
        RECT 0.425000 1.495000 3.070000 1.665000 ;
        RECT 2.415000 1.415000 3.070000 1.495000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.285000 0.255000 3.615000 0.905000 ;
        RECT 3.285000 1.495000 3.615000 2.465000 ;
        RECT 3.445000 0.905000 3.615000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.280000 0.525000 0.655000 ;
      RECT 0.085000  0.655000 3.105000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.835000 ;
      RECT 0.085000  1.835000 2.085000 2.005000 ;
      RECT 0.085000  2.005000 0.615000 2.465000 ;
      RECT 0.975000  0.085000 1.305000 0.485000 ;
      RECT 0.975000  2.175000 1.305000 2.635000 ;
      RECT 1.755000  0.255000 2.085000 0.655000 ;
      RECT 1.755000  2.005000 2.085000 2.465000 ;
      RECT 2.535000  1.835000 2.860000 2.635000 ;
      RECT 2.635000  0.085000 2.965000 0.485000 ;
      RECT 2.925000  0.825000 3.105000 1.075000 ;
      RECT 2.925000  1.075000 3.275000 1.245000 ;
      RECT 3.785000  0.085000 4.055000 0.905000 ;
      RECT 3.785000  1.495000 4.055000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__maj3_2
MACRO sky130_fd_sc_hd__maj3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__maj3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 1.075000 1.450000 1.635000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.960000 1.075000 2.290000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 0.890000 1.285000 ;
        RECT 0.720000 1.285000 0.890000 1.915000 ;
        RECT 0.720000 1.915000 1.790000 2.085000 ;
        RECT 1.620000 2.085000 1.790000 2.225000 ;
        RECT 1.620000 2.225000 2.630000 2.395000 ;
        RECT 2.460000 1.075000 2.945000 1.245000 ;
        RECT 2.460000 1.245000 2.630000 2.225000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.375000 0.255000 3.705000 0.490000 ;
        RECT 3.375000 1.455000 4.975000 1.625000 ;
        RECT 3.375000 1.625000 3.705000 2.465000 ;
        RECT 3.455000 0.490000 3.705000 0.715000 ;
        RECT 3.455000 0.715000 4.975000 0.905000 ;
        RECT 4.215000 0.255000 4.545000 0.715000 ;
        RECT 4.215000 1.625000 4.545000 2.465000 ;
        RECT 4.715000 0.905000 4.975000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.085000 0.310000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.255000 0.635000 0.660000 ;
      RECT 0.085000  0.660000 2.290000 0.715000 ;
      RECT 0.085000  0.715000 3.285000 0.885000 ;
      RECT 0.085000  0.885000 0.255000 1.455000 ;
      RECT 0.085000  1.455000 0.465000 2.465000 ;
      RECT 1.120000  0.085000 1.450000 0.490000 ;
      RECT 1.120000  2.255000 1.450000 2.635000 ;
      RECT 1.620000  0.885000 1.790000 1.545000 ;
      RECT 1.620000  1.545000 2.290000 1.745000 ;
      RECT 1.960000  0.255000 2.290000 0.660000 ;
      RECT 1.960000  1.745000 2.290000 2.055000 ;
      RECT 2.845000  1.455000 3.175000 2.635000 ;
      RECT 2.860000  0.085000 3.205000 0.545000 ;
      RECT 3.115000  0.885000 3.285000 1.075000 ;
      RECT 3.115000  1.075000 4.545000 1.285000 ;
      RECT 3.875000  0.085000 4.045000 0.545000 ;
      RECT 3.875000  1.795000 4.045000 2.635000 ;
      RECT 4.715000  0.085000 4.885000 0.545000 ;
      RECT 4.715000  1.795000 4.925000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__maj3_4
MACRO sky130_fd_sc_hd__mux2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 0.255000 2.265000 1.415000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.615000 0.815000 1.785000 1.615000 ;
        RECT 1.615000 1.615000 2.625000 1.785000 ;
        RECT 2.435000 0.255000 2.625000 1.615000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.910000 0.995000 1.105000 1.325000 ;
        RECT 0.935000 1.325000 1.105000 2.295000 ;
        RECT 0.935000 2.295000 2.965000 2.465000 ;
        RECT 2.795000 1.440000 3.545000 1.630000 ;
        RECT 2.795000 1.630000 2.965000 2.295000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.255000 0.345000 0.825000 ;
        RECT 0.090000 0.825000 0.260000 1.495000 ;
        RECT 0.090000 1.495000 0.425000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.420000 -0.085000 0.590000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.430000  0.995000 0.685000 1.325000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 0.515000  0.655000 1.445000 0.825000 ;
      RECT 0.515000  0.825000 0.685000 0.995000 ;
      RECT 0.595000  1.495000 0.765000 2.635000 ;
      RECT 1.270000  0.255000 1.800000 0.620000 ;
      RECT 1.270000  0.620000 1.445000 0.655000 ;
      RECT 1.275000  0.825000 1.445000 1.955000 ;
      RECT 1.275000  1.955000 2.400000 2.125000 ;
      RECT 2.805000  0.085000 3.315000 0.620000 ;
      RECT 2.825000  0.895000 4.055000 1.065000 ;
      RECT 3.135000  1.875000 3.305000 2.635000 ;
      RECT 3.535000  0.290000 3.780000 0.895000 ;
      RECT 3.540000  1.875000 4.055000 2.285000 ;
      RECT 3.715000  1.065000 4.055000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__mux2_1
MACRO sky130_fd_sc_hd__mux2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.815000 0.765000 2.445000 1.280000 ;
        RECT 2.275000 1.280000 2.445000 1.315000 ;
        RECT 2.275000 1.315000 3.090000 1.625000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.625000 0.735000 3.090000 1.025000 ;
        RECT 2.900000 0.420000 3.090000 0.735000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.360000 0.755000 3.550000 1.625000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.765000 0.750000 ;
        RECT 0.515000 0.750000 0.685000 1.595000 ;
        RECT 0.515000 1.595000 0.825000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.085000 0.345000 0.885000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.855000  0.995000 1.165000 1.325000 ;
      RECT 0.935000  0.085000 1.265000 0.465000 ;
      RECT 0.995000  0.635000 1.605000 0.805000 ;
      RECT 0.995000  0.805000 1.165000 0.995000 ;
      RECT 0.995000  1.325000 1.165000 1.835000 ;
      RECT 0.995000  1.835000 1.655000 2.005000 ;
      RECT 1.025000  2.175000 1.315000 2.635000 ;
      RECT 1.335000  0.995000 1.505000 1.495000 ;
      RECT 1.335000  1.495000 1.995000 1.665000 ;
      RECT 1.435000  0.295000 2.730000 0.465000 ;
      RECT 1.435000  0.465000 1.605000 0.635000 ;
      RECT 1.485000  2.005000 1.655000 2.255000 ;
      RECT 1.485000  2.255000 2.795000 2.425000 ;
      RECT 1.825000  1.665000 1.995000 1.835000 ;
      RECT 1.825000  1.835000 4.050000 2.005000 ;
      RECT 3.325000  2.175000 3.545000 2.635000 ;
      RECT 3.350000  0.085000 3.550000 0.585000 ;
      RECT 3.715000  2.005000 4.050000 2.465000 ;
      RECT 3.720000  0.255000 4.050000 1.835000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__mux2_2
MACRO sky130_fd_sc_hd__mux2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 0.995000 1.750000 1.615000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 0.995000 2.435000 1.325000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.995000 0.740000 1.325000 ;
        RECT 0.570000 0.635000 2.850000 0.805000 ;
        RECT 0.570000 0.805000 0.740000 0.995000 ;
        RECT 2.680000 0.805000 2.850000 0.995000 ;
        RECT 2.680000 0.995000 3.395000 1.325000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.915000 0.255000 4.085000 0.635000 ;
        RECT 3.915000 0.635000 5.430000 0.805000 ;
        RECT 3.915000 1.575000 5.430000 1.745000 ;
        RECT 3.915000 1.745000 4.085000 2.465000 ;
        RECT 4.755000 0.255000 4.925000 0.635000 ;
        RECT 4.755000 1.745000 4.925000 2.465000 ;
        RECT 5.200000 0.805000 5.430000 1.575000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.090000  0.295000 0.345000 0.625000 ;
      RECT 0.090000  0.625000 0.260000 1.495000 ;
      RECT 0.090000  1.495000 1.080000 1.665000 ;
      RECT 0.090000  1.665000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  1.835000 0.820000 2.635000 ;
      RECT 0.910000  0.995000 1.080000 1.495000 ;
      RECT 0.990000  1.935000 1.340000 2.275000 ;
      RECT 0.990000  2.275000 2.770000 2.445000 ;
      RECT 1.530000  1.935000 3.245000 2.105000 ;
      RECT 1.975000  0.295000 3.230000 0.465000 ;
      RECT 1.980000  1.595000 3.735000 1.765000 ;
      RECT 3.060000  0.465000 3.230000 0.655000 ;
      RECT 3.060000  0.655000 3.735000 0.825000 ;
      RECT 3.075000  2.105000 3.245000 2.465000 ;
      RECT 3.415000  0.085000 3.745000 0.465000 ;
      RECT 3.415000  2.255000 3.745000 2.635000 ;
      RECT 3.565000  0.825000 3.735000 1.075000 ;
      RECT 3.565000  1.075000 5.030000 1.245000 ;
      RECT 3.565000  1.245000 3.735000 1.595000 ;
      RECT 3.565000  1.765000 3.735000 1.785000 ;
      RECT 4.255000  0.085000 4.585000 0.465000 ;
      RECT 4.255000  1.915000 4.585000 2.635000 ;
      RECT 5.095000  0.085000 5.425000 0.465000 ;
      RECT 5.095000  1.915000 5.425000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__mux2_4
MACRO sky130_fd_sc_hd__mux2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.180000 0.645000 6.895000 0.815000 ;
        RECT 5.180000 0.815000 5.350000 1.325000 ;
        RECT 5.305000 0.425000 5.890000 0.645000 ;
        RECT 6.725000 0.815000 6.895000 0.995000 ;
        RECT 6.725000 0.995000 7.195000 1.165000 ;
        RECT 7.025000 1.165000 7.195000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.290000 1.105000 4.475000 1.275000 ;
        RECT 4.305000 0.995000 4.475000 1.105000 ;
        RECT 4.305000 1.275000 4.475000 1.325000 ;
      LAYER mcon ;
        RECT 4.290000 1.105000 4.460000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.960000 0.995000 8.245000 1.325000 ;
      LAYER mcon ;
        RECT 7.960000 1.105000 8.130000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.230000 1.075000 4.520000 1.120000 ;
        RECT 4.230000 1.120000 8.190000 1.260000 ;
        RECT 4.230000 1.260000 4.520000 1.305000 ;
        RECT 7.900000 1.075000 8.190000 1.120000 ;
        RECT 7.900000 1.260000 8.190000 1.305000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.739500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.795000 0.995000 3.965000 1.495000 ;
        RECT 3.795000 1.495000 6.035000 1.665000 ;
        RECT 5.670000 0.995000 6.035000 1.495000 ;
      LAYER mcon ;
        RECT 5.670000 1.445000 5.840000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.215000 0.995000 9.510000 1.615000 ;
      LAYER mcon ;
        RECT 9.340000 1.445000 9.510000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.610000 1.415000 5.900000 1.460000 ;
        RECT 5.610000 1.460000 9.570000 1.600000 ;
        RECT 5.610000 1.600000 5.900000 1.645000 ;
        RECT 9.280000 1.415000 9.570000 1.460000 ;
        RECT 9.280000 1.600000 9.570000 1.645000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.255000 0.765000 0.635000 ;
        RECT 0.595000 0.635000 3.285000 0.805000 ;
        RECT 0.595000 0.805000 0.815000 1.575000 ;
        RECT 0.595000 1.575000 3.285000 1.745000 ;
        RECT 0.595000 1.745000 0.765000 2.465000 ;
        RECT 1.435000 0.295000 1.605000 0.635000 ;
        RECT 1.435000 1.745000 1.605000 2.465000 ;
        RECT 2.275000 0.255000 2.445000 0.635000 ;
        RECT 2.275000 1.745000 2.445000 2.465000 ;
        RECT 3.115000 0.295000 3.285000 0.635000 ;
        RECT 3.115000 1.745000 3.285000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.465000 ;
      RECT 0.090000  1.915000 0.425000 2.635000 ;
      RECT 0.935000  0.085000 1.265000 0.465000 ;
      RECT 0.935000  1.915000 1.265000 2.635000 ;
      RECT 0.985000  1.075000 3.625000 1.245000 ;
      RECT 1.775000  0.085000 2.105000 0.465000 ;
      RECT 1.775000  1.915000 2.105000 2.635000 ;
      RECT 2.615000  0.085000 2.945000 0.465000 ;
      RECT 2.615000  1.915000 2.945000 2.635000 ;
      RECT 3.455000  0.085000 3.785000 0.465000 ;
      RECT 3.455000  0.635000 4.920000 0.805000 ;
      RECT 3.455000  0.805000 3.625000 1.075000 ;
      RECT 3.455000  1.245000 3.625000 1.835000 ;
      RECT 3.455000  1.835000 8.225000 2.005000 ;
      RECT 3.455000  2.255000 3.785000 2.635000 ;
      RECT 3.955000  0.295000 5.125000 0.465000 ;
      RECT 3.955000  2.255000 5.905000 2.425000 ;
      RECT 4.750000  0.805000 4.920000 0.935000 ;
      RECT 6.060000  0.085000 6.390000 0.465000 ;
      RECT 6.075000  2.175000 6.245000 2.635000 ;
      RECT 6.345000  0.995000 6.515000 1.495000 ;
      RECT 6.345000  1.495000 8.855000 1.665000 ;
      RECT 6.480000  2.255000 8.645000 2.425000 ;
      RECT 6.575000  0.295000 7.865000 0.465000 ;
      RECT 7.115000  0.635000 7.670000 0.805000 ;
      RECT 7.500000  0.805000 7.670000 0.935000 ;
      RECT 8.685000  0.645000 9.485000 0.815000 ;
      RECT 8.685000  0.815000 8.855000 1.495000 ;
      RECT 8.685000  1.665000 8.855000 1.915000 ;
      RECT 8.685000  1.915000 9.485000 2.085000 ;
      RECT 8.815000  0.085000 9.145000 0.465000 ;
      RECT 8.815000  2.255000 9.145000 2.635000 ;
      RECT 9.315000  0.295000 9.485000 0.645000 ;
      RECT 9.315000  1.795000 9.485000 1.915000 ;
      RECT 9.315000  2.085000 9.485000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 4.750000  0.765000 4.920000 0.935000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.500000  0.765000 7.670000 0.935000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 4.690000 0.735000 4.980000 0.780000 ;
      RECT 4.690000 0.780000 7.730000 0.920000 ;
      RECT 4.690000 0.920000 4.980000 0.965000 ;
      RECT 7.440000 0.735000 7.730000 0.780000 ;
      RECT 7.440000 0.920000 7.730000 0.965000 ;
  END
END sky130_fd_sc_hd__mux2_8
MACRO sky130_fd_sc_hd__mux2i_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2i_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.060000 0.420000 1.285000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 0.995000 1.125000 1.155000 ;
        RECT 0.955000 1.155000 1.205000 1.325000 ;
        RECT 1.035000 1.325000 1.205000 1.445000 ;
        RECT 1.035000 1.445000 1.235000 2.110000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.260000 0.760000 3.595000 1.620000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  0.480500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.590000 0.595000 0.780000 1.455000 ;
        RECT 0.590000 1.455000 0.840000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.255000 1.805000 0.425000 ;
      RECT 0.085000  0.425000 0.440000 0.465000 ;
      RECT 0.085000  0.465000 0.345000 0.885000 ;
      RECT 0.120000  1.455000 0.420000 2.295000 ;
      RECT 0.120000  2.295000 1.575000 2.465000 ;
      RECT 0.955000  0.655000 1.520000 0.715000 ;
      RECT 0.955000  0.715000 2.620000 0.825000 ;
      RECT 0.965000  0.425000 1.805000 0.465000 ;
      RECT 1.295000  0.825000 2.620000 0.885000 ;
      RECT 1.385000  1.075000 3.085000 1.310000 ;
      RECT 1.405000  1.480000 2.615000 1.650000 ;
      RECT 1.405000  1.650000 1.575000 2.295000 ;
      RECT 1.745000  1.835000 1.975000 2.635000 ;
      RECT 1.975000  0.085000 2.145000 0.545000 ;
      RECT 2.285000  1.650000 2.615000 2.465000 ;
      RECT 2.385000  0.255000 2.620000 0.715000 ;
      RECT 2.800000  0.255000 3.165000 0.485000 ;
      RECT 2.800000  0.485000 3.085000 1.075000 ;
      RECT 2.860000  1.310000 3.085000 2.465000 ;
      RECT 3.295000  1.835000 3.590000 2.635000 ;
      RECT 3.335000  0.085000 3.555000 0.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__mux2i_1
MACRO sky130_fd_sc_hd__mux2i_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2i_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.470000 1.075000 3.560000 1.275000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.310000 0.995000 4.635000 1.615000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.995000 0.780000 1.325000 ;
        RECT 0.580000 0.725000 0.780000 0.995000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  1.691250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.715000 0.295000 4.975000 0.465000 ;
        RECT 2.715000 2.255000 4.975000 2.425000 ;
        RECT 4.750000 1.785000 4.975000 2.255000 ;
        RECT 4.805000 0.465000 4.975000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.675000 ;
      RECT 0.085000  0.675000 0.260000 1.495000 ;
      RECT 0.085000  1.495000 1.395000 1.665000 ;
      RECT 0.085000  1.665000 0.260000 2.135000 ;
      RECT 0.085000  2.135000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.835000 0.545000 ;
      RECT 0.515000  2.255000 0.845000 2.635000 ;
      RECT 0.935000  1.835000 1.735000 2.005000 ;
      RECT 1.015000  0.575000 1.255000 0.935000 ;
      RECT 1.225000  1.155000 1.985000 1.325000 ;
      RECT 1.225000  1.325000 1.395000 1.495000 ;
      RECT 1.355000  2.255000 1.685000 2.635000 ;
      RECT 1.435000  0.085000 1.685000 0.885000 ;
      RECT 1.565000  1.495000 3.465000 1.665000 ;
      RECT 1.565000  1.665000 1.735000 1.835000 ;
      RECT 1.655000  1.075000 1.985000 1.155000 ;
      RECT 1.855000  0.295000 2.025000 0.735000 ;
      RECT 1.855000  0.735000 3.465000 0.905000 ;
      RECT 1.855000  2.135000 2.080000 2.465000 ;
      RECT 1.910000  1.835000 2.885000 1.915000 ;
      RECT 1.910000  1.915000 4.350000 2.005000 ;
      RECT 1.910000  2.005000 2.080000 2.135000 ;
      RECT 2.275000  0.085000 2.445000 0.545000 ;
      RECT 2.275000  2.175000 2.525000 2.635000 ;
      RECT 2.715000  2.005000 4.350000 2.085000 ;
      RECT 3.135000  0.655000 3.465000 0.735000 ;
      RECT 3.135000  1.665000 3.465000 1.715000 ;
      RECT 3.850000  0.655000 4.345000 0.825000 ;
      RECT 3.850000  0.825000 4.105000 0.935000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  0.765000 1.240000 0.935000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 3.850000  0.765000 4.020000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
    LAYER met1 ;
      RECT 1.010000 0.735000 1.300000 0.780000 ;
      RECT 1.010000 0.780000 4.080000 0.920000 ;
      RECT 1.010000 0.920000 1.300000 0.965000 ;
      RECT 3.790000 0.735000 4.080000 0.780000 ;
      RECT 3.790000 0.920000 4.080000 0.965000 ;
  END
END sky130_fd_sc_hd__mux2i_2
MACRO sky130_fd_sc_hd__mux2i_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2i_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 0.995000 1.070000 1.105000 ;
        RECT 0.560000 1.105000 1.240000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 0.995000 3.550000 1.325000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  1.237500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.845000 1.075000 5.930000 1.290000 ;
        RECT 5.760000 1.290000 5.930000 1.425000 ;
        RECT 5.760000 1.425000 7.850000 1.595000 ;
        RECT 7.680000 0.995000 7.850000 1.425000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  2.194500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.315000 3.785000 0.485000 ;
        RECT 0.095000 0.485000 0.320000 2.255000 ;
        RECT 0.095000 2.255000 3.785000 2.425000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.515000  0.655000 1.700000 0.825000 ;
      RECT 0.515000  1.575000 5.580000 1.745000 ;
      RECT 1.355000  0.825000 1.700000 0.935000 ;
      RECT 2.195000  0.655000 5.485000 0.825000 ;
      RECT 2.195000  1.915000 7.165000 2.085000 ;
      RECT 3.975000  0.085000 4.305000 0.465000 ;
      RECT 3.975000  2.255000 4.305000 2.635000 ;
      RECT 4.475000  0.255000 4.645000 0.655000 ;
      RECT 4.815000  0.085000 5.145000 0.465000 ;
      RECT 4.815000  2.255000 5.145000 2.635000 ;
      RECT 5.315000  0.255000 5.485000 0.655000 ;
      RECT 5.655000  0.085000 5.980000 0.590000 ;
      RECT 5.655000  2.255000 5.985000 2.635000 ;
      RECT 6.150000  0.255000 6.325000 0.715000 ;
      RECT 6.150000  0.715000 7.165000 0.905000 ;
      RECT 6.150000  0.905000 6.450000 0.935000 ;
      RECT 6.155000  1.795000 6.325000 1.915000 ;
      RECT 6.155000  2.085000 6.325000 2.465000 ;
      RECT 6.495000  2.255000 6.825000 2.635000 ;
      RECT 6.545000  0.085000 6.795000 0.545000 ;
      RECT 6.730000  1.075000 7.510000 1.245000 ;
      RECT 6.995000  0.510000 7.165000 0.715000 ;
      RECT 6.995000  1.795000 7.165000 1.915000 ;
      RECT 6.995000  2.085000 7.165000 2.465000 ;
      RECT 7.340000  0.655000 8.195000 0.825000 ;
      RECT 7.340000  0.825000 7.510000 1.075000 ;
      RECT 7.435000  0.085000 7.765000 0.465000 ;
      RECT 7.435000  2.255000 7.765000 2.635000 ;
      RECT 7.935000  0.255000 8.195000 0.655000 ;
      RECT 7.935000  1.795000 8.195000 2.465000 ;
      RECT 8.020000  0.825000 8.195000 1.795000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.530000  0.765000 1.700000 0.935000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.150000  0.765000 6.320000 0.935000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
    LAYER met1 ;
      RECT 1.470000 0.735000 1.760000 0.780000 ;
      RECT 1.470000 0.780000 6.380000 0.920000 ;
      RECT 1.470000 0.920000 1.760000 0.965000 ;
      RECT 6.090000 0.735000 6.380000 0.780000 ;
      RECT 6.090000 0.920000 6.380000 0.965000 ;
  END
END sky130_fd_sc_hd__mux2i_4
MACRO sky130_fd_sc_hd__mux4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 0.995000 1.240000 1.615000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.995000 0.495000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.250000 1.055000 5.580000 1.675000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.800000 1.055000 5.045000 1.675000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.265000 0.995000 3.565000 1.995000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.055000 0.995000 6.345000 1.675000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.315000 0.255000 9.575000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.175000  0.260000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 1.185000 0.805000 ;
      RECT 0.175000  1.795000 1.705000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.255000 0.845000 2.635000 ;
      RECT 1.015000  0.255000 2.090000 0.425000 ;
      RECT 1.015000  0.425000 1.185000 0.635000 ;
      RECT 1.015000  2.135000 1.185000 2.295000 ;
      RECT 1.015000  2.295000 2.545000 2.465000 ;
      RECT 1.410000  0.595000 1.750000 0.765000 ;
      RECT 1.410000  0.765000 1.700000 0.935000 ;
      RECT 1.410000  0.935000 1.580000 1.455000 ;
      RECT 1.410000  1.455000 2.045000 1.625000 ;
      RECT 1.535000  1.965000 1.705000 2.125000 ;
      RECT 1.875000  1.625000 2.045000 1.955000 ;
      RECT 1.875000  1.955000 2.205000 2.125000 ;
      RECT 1.920000  0.425000 2.090000 0.760000 ;
      RECT 2.080000  1.105000 2.620000 1.285000 ;
      RECT 2.260000  0.430000 2.620000 1.105000 ;
      RECT 2.260000  1.285000 2.620000 1.395000 ;
      RECT 2.260000  1.395000 3.065000 1.625000 ;
      RECT 2.375000  1.795000 2.545000 2.295000 ;
      RECT 2.715000  1.625000 3.065000 2.465000 ;
      RECT 2.800000  0.085000 3.090000 0.805000 ;
      RECT 3.235000  2.255000 3.565000 2.635000 ;
      RECT 3.380000  0.255000 4.980000 0.425000 ;
      RECT 3.380000  0.425000 3.550000 0.795000 ;
      RECT 3.720000  0.595000 4.050000 0.845000 ;
      RECT 3.735000  0.845000 4.050000 0.920000 ;
      RECT 3.735000  0.920000 3.905000 1.445000 ;
      RECT 3.735000  1.445000 4.495000 1.615000 ;
      RECT 3.825000  1.785000 3.995000 2.295000 ;
      RECT 3.825000  2.295000 4.835000 2.465000 ;
      RECT 4.075000  1.095000 4.405000 1.105000 ;
      RECT 4.075000  1.105000 4.460000 1.265000 ;
      RECT 4.165000  1.615000 4.495000 2.125000 ;
      RECT 4.220000  0.595000 4.390000 0.715000 ;
      RECT 4.220000  0.715000 5.740000 0.885000 ;
      RECT 4.220000  0.885000 4.390000 0.925000 ;
      RECT 4.290000  1.265000 4.460000 1.275000 ;
      RECT 4.625000  0.425000 4.980000 0.465000 ;
      RECT 4.665000  1.915000 5.730000 2.085000 ;
      RECT 4.665000  2.085000 4.835000 2.295000 ;
      RECT 5.060000  2.255000 5.390000 2.635000 ;
      RECT 5.150000  0.085000 5.320000 0.545000 ;
      RECT 5.495000  0.295000 5.740000 0.715000 ;
      RECT 5.560000  2.085000 5.730000 2.465000 ;
      RECT 5.980000  2.255000 6.330000 2.635000 ;
      RECT 6.010000  0.085000 6.340000 0.465000 ;
      RECT 6.500000  2.135000 6.685000 2.465000 ;
      RECT 6.510000  0.325000 6.685000 0.655000 ;
      RECT 6.515000  0.655000 6.685000 1.105000 ;
      RECT 6.515000  1.105000 6.805000 1.275000 ;
      RECT 6.515000  1.275000 6.685000 2.135000 ;
      RECT 6.980000  0.765000 7.220000 0.935000 ;
      RECT 6.980000  0.935000 7.150000 2.135000 ;
      RECT 6.980000  2.135000 7.190000 2.465000 ;
      RECT 7.030000  0.255000 7.200000 0.415000 ;
      RECT 7.030000  0.415000 7.560000 0.585000 ;
      RECT 7.360000  2.255000 7.690000 2.295000 ;
      RECT 7.360000  2.295000 8.645000 2.465000 ;
      RECT 7.390000  0.585000 7.560000 1.755000 ;
      RECT 7.390000  1.755000 8.175000 1.985000 ;
      RECT 7.730000  0.255000 8.725000 0.425000 ;
      RECT 7.730000  0.425000 7.900000 0.585000 ;
      RECT 7.845000  1.985000 8.175000 2.125000 ;
      RECT 7.970000  0.765000 8.385000 0.925000 ;
      RECT 7.970000  0.925000 8.380000 0.935000 ;
      RECT 8.190000  1.105000 8.645000 1.275000 ;
      RECT 8.210000  0.595000 8.385000 0.765000 ;
      RECT 8.475000  1.665000 9.125000 1.835000 ;
      RECT 8.475000  1.835000 8.645000 2.295000 ;
      RECT 8.555000  0.425000 8.725000 0.715000 ;
      RECT 8.555000  0.715000 9.125000 0.885000 ;
      RECT 8.815000  2.255000 9.145000 2.635000 ;
      RECT 8.895000  0.085000 9.065000 0.545000 ;
      RECT 8.955000  0.885000 9.125000 1.665000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.530000  0.765000 1.700000 0.935000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.450000  1.105000 2.620000 1.275000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.290000  1.105000 4.460000 1.275000 ;
      RECT 4.325000  1.785000 4.495000 1.955000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.635000  1.105000 6.805000 1.275000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.050000  0.765000 7.220000 0.935000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.555000  1.785000 7.725000 1.955000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.475000  1.105000 8.645000 1.275000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 1.470000 0.735000 1.760000 0.780000 ;
      RECT 1.470000 0.780000 8.200000 0.920000 ;
      RECT 1.470000 0.920000 1.760000 0.965000 ;
      RECT 2.390000 1.075000 2.680000 1.120000 ;
      RECT 2.390000 1.120000 4.520000 1.260000 ;
      RECT 2.390000 1.260000 2.680000 1.305000 ;
      RECT 4.230000 1.075000 4.520000 1.120000 ;
      RECT 4.230000 1.260000 4.520000 1.305000 ;
      RECT 4.265000 1.755000 4.555000 1.800000 ;
      RECT 4.265000 1.800000 7.785000 1.940000 ;
      RECT 4.265000 1.940000 4.555000 1.985000 ;
      RECT 6.575000 1.075000 6.865000 1.120000 ;
      RECT 6.575000 1.120000 8.705000 1.260000 ;
      RECT 6.575000 1.260000 6.865000 1.305000 ;
      RECT 6.990000 0.735000 7.280000 0.780000 ;
      RECT 6.990000 0.920000 7.280000 0.965000 ;
      RECT 7.495000 1.755000 7.785000 1.800000 ;
      RECT 7.495000 1.940000 7.785000 1.985000 ;
      RECT 7.910000 0.735000 8.200000 0.780000 ;
      RECT 7.910000 0.920000 8.200000 0.965000 ;
      RECT 8.415000 1.075000 8.705000 1.120000 ;
      RECT 8.415000 1.260000 8.705000 1.305000 ;
  END
END sky130_fd_sc_hd__mux4_1
MACRO sky130_fd_sc_hd__mux4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.535000 0.375000 6.845000 0.995000 ;
        RECT 6.535000 0.995000 6.945000 1.075000 ;
        RECT 6.635000 1.075000 6.945000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.745000 0.715000 5.115000 1.395000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835000 0.765000 1.235000 1.095000 ;
        RECT 1.020000 0.395000 1.235000 0.765000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.240000 0.715000 2.615000 1.015000 ;
        RECT 2.410000 1.015000 2.615000 1.320000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.393000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.975000 0.325000 1.745000 ;
      LAYER mcon ;
        RECT 0.145000 1.445000 0.315000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.005000 1.445000 1.390000 1.615000 ;
        RECT 1.220000 1.285000 1.390000 1.445000 ;
      LAYER mcon ;
        RECT 1.065000 1.445000 1.235000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.125000 1.245000 6.465000 1.645000 ;
      LAYER mcon ;
        RECT 6.125000 1.445000 6.295000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.085000 1.415000 0.375000 1.460000 ;
        RECT 0.085000 1.460000 6.355000 1.600000 ;
        RECT 0.085000 1.600000 0.375000 1.645000 ;
        RECT 1.005000 1.415000 1.295000 1.460000 ;
        RECT 1.005000 1.600000 1.295000 1.645000 ;
        RECT 6.065000 1.415000 6.355000 1.460000 ;
        RECT 6.065000 1.600000 6.355000 1.645000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.303000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 0.715000 3.075000 1.320000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.355000 1.835000 7.765000 2.455000 ;
        RECT 7.435000 0.265000 7.765000 0.725000 ;
        RECT 7.455000 1.495000 7.765000 1.835000 ;
        RECT 7.595000 0.725000 7.765000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.170000  0.345000 0.345000 0.635000 ;
      RECT 0.170000  0.635000 0.665000 0.805000 ;
      RECT 0.175000  1.915000 1.900000 1.955000 ;
      RECT 0.175000  1.955000 0.665000 2.085000 ;
      RECT 0.175000  2.085000 0.345000 2.375000 ;
      RECT 0.495000  0.805000 0.665000 1.785000 ;
      RECT 0.495000  1.785000 1.900000 1.915000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.255000 0.845000 2.635000 ;
      RECT 1.405000  0.705000 1.730000 1.035000 ;
      RECT 1.410000  2.125000 2.240000 2.295000 ;
      RECT 1.470000  0.365000 2.070000 0.535000 ;
      RECT 1.560000  1.035000 1.730000 1.575000 ;
      RECT 1.560000  1.575000 1.900000 1.785000 ;
      RECT 1.900000  0.535000 2.070000 1.235000 ;
      RECT 1.900000  1.235000 2.240000 1.405000 ;
      RECT 2.070000  1.405000 2.240000 2.125000 ;
      RECT 2.450000  0.085000 2.780000 0.545000 ;
      RECT 2.595000  2.055000 2.825000 2.635000 ;
      RECT 2.970000  1.785000 3.315000 1.955000 ;
      RECT 2.985000  0.295000 3.415000 0.465000 ;
      RECT 3.145000  1.490000 3.415000 1.660000 ;
      RECT 3.145000  1.660000 3.315000 1.785000 ;
      RECT 3.245000  0.465000 3.415000 1.060000 ;
      RECT 3.245000  1.060000 3.480000 1.390000 ;
      RECT 3.245000  1.390000 3.415000 1.490000 ;
      RECT 3.305000  2.125000 3.820000 2.295000 ;
      RECT 3.565000  1.810000 3.820000 2.125000 ;
      RECT 3.585000  0.345000 3.820000 0.675000 ;
      RECT 3.650000  0.675000 3.820000 1.810000 ;
      RECT 3.990000  0.345000 4.180000 2.125000 ;
      RECT 3.990000  2.125000 4.515000 2.295000 ;
      RECT 4.395000  0.255000 4.600000 0.585000 ;
      RECT 4.395000  0.585000 4.565000 1.565000 ;
      RECT 4.395000  1.565000 5.495000 1.735000 ;
      RECT 4.395000  1.735000 4.585000 1.895000 ;
      RECT 4.755000  2.005000 5.100000 2.635000 ;
      RECT 4.795000  0.085000 5.125000 0.545000 ;
      RECT 5.325000  0.295000 6.220000 0.465000 ;
      RECT 5.325000  0.465000 5.495000 1.565000 ;
      RECT 5.325000  1.735000 5.495000 2.155000 ;
      RECT 5.325000  2.155000 6.275000 2.325000 ;
      RECT 5.665000  0.705000 6.285000 1.035000 ;
      RECT 5.665000  1.035000 5.955000 1.985000 ;
      RECT 6.525000  2.125000 6.845000 2.295000 ;
      RECT 6.675000  1.495000 7.285000 1.665000 ;
      RECT 6.675000  1.665000 6.845000 2.125000 ;
      RECT 7.015000  0.085000 7.265000 0.815000 ;
      RECT 7.015000  1.835000 7.185000 2.635000 ;
      RECT 7.115000  0.995000 7.425000 1.325000 ;
      RECT 7.115000  1.325000 7.285000 1.495000 ;
      RECT 7.935000  0.085000 8.190000 0.885000 ;
      RECT 7.935000  1.495000 8.185000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  1.785000 1.695000 1.955000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.125000 2.155000 2.295000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.125000 3.535000 2.295000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.125000 4.455000 2.295000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  1.785000 5.835000 1.955000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.125000 6.755000 2.295000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
    LAYER met1 ;
      RECT 1.465000 1.755000 1.755000 1.800000 ;
      RECT 1.465000 1.800000 5.895000 1.940000 ;
      RECT 1.465000 1.940000 1.755000 1.985000 ;
      RECT 1.925000 2.095000 2.215000 2.140000 ;
      RECT 1.925000 2.140000 3.595000 2.280000 ;
      RECT 1.925000 2.280000 2.215000 2.325000 ;
      RECT 3.305000 2.095000 3.595000 2.140000 ;
      RECT 3.305000 2.280000 3.595000 2.325000 ;
      RECT 4.225000 2.095000 4.515000 2.140000 ;
      RECT 4.225000 2.140000 6.815000 2.280000 ;
      RECT 4.225000 2.280000 4.515000 2.325000 ;
      RECT 5.605000 1.755000 5.895000 1.800000 ;
      RECT 5.605000 1.940000 5.895000 1.985000 ;
      RECT 6.525000 2.095000 6.815000 2.140000 ;
      RECT 6.525000 2.280000 6.815000 2.325000 ;
  END
END sky130_fd_sc_hd__mux4_2
MACRO sky130_fd_sc_hd__mux4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.540000 0.375000 6.850000 0.995000 ;
        RECT 6.540000 0.995000 6.950000 1.075000 ;
        RECT 6.640000 1.075000 6.950000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.750000 0.715000 5.120000 1.395000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.840000 0.765000 1.240000 1.095000 ;
        RECT 1.025000 0.395000 1.240000 0.765000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.245000 0.715000 2.620000 1.015000 ;
        RECT 2.415000 1.015000 2.620000 1.320000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.393000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.975000 0.330000 1.745000 ;
      LAYER mcon ;
        RECT 0.150000 1.445000 0.320000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.010000 1.445000 1.395000 1.615000 ;
        RECT 1.225000 1.285000 1.395000 1.445000 ;
      LAYER mcon ;
        RECT 1.070000 1.445000 1.240000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.130000 1.245000 6.470000 1.645000 ;
      LAYER mcon ;
        RECT 6.130000 1.445000 6.300000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.085000 1.415000 0.380000 1.460000 ;
        RECT 0.085000 1.460000 6.360000 1.600000 ;
        RECT 0.085000 1.600000 0.380000 1.645000 ;
        RECT 1.010000 1.415000 1.300000 1.460000 ;
        RECT 1.010000 1.600000 1.300000 1.645000 ;
        RECT 6.070000 1.415000 6.360000 1.460000 ;
        RECT 6.070000 1.600000 6.360000 1.645000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.303000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 0.715000 3.080000 1.320000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.360000 1.835000 7.770000 2.455000 ;
        RECT 7.440000 0.265000 7.770000 0.725000 ;
        RECT 7.460000 1.495000 7.770000 1.835000 ;
        RECT 7.600000 0.725000 7.770000 1.065000 ;
        RECT 7.600000 1.065000 8.685000 1.305000 ;
        RECT 7.600000 1.305000 7.770000 1.495000 ;
        RECT 8.360000 0.265000 8.685000 1.065000 ;
        RECT 8.360000 1.305000 8.685000 2.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.135000  0.345000 0.345000 0.635000 ;
      RECT 0.135000  0.635000 0.670000 0.805000 ;
      RECT 0.135000  1.915000 1.905000 1.955000 ;
      RECT 0.135000  1.955000 0.670000 2.085000 ;
      RECT 0.135000  2.085000 0.345000 2.375000 ;
      RECT 0.500000  0.805000 0.670000 1.785000 ;
      RECT 0.500000  1.785000 1.905000 1.915000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.255000 0.845000 2.635000 ;
      RECT 1.410000  0.705000 1.735000 1.035000 ;
      RECT 1.415000  2.125000 2.245000 2.295000 ;
      RECT 1.475000  0.365000 2.075000 0.535000 ;
      RECT 1.565000  1.035000 1.735000 1.575000 ;
      RECT 1.565000  1.575000 1.905000 1.785000 ;
      RECT 1.905000  0.535000 2.075000 1.235000 ;
      RECT 1.905000  1.235000 2.245000 1.405000 ;
      RECT 2.075000  1.405000 2.245000 2.125000 ;
      RECT 2.455000  0.085000 2.785000 0.545000 ;
      RECT 2.600000  2.055000 2.830000 2.635000 ;
      RECT 2.975000  1.785000 3.320000 1.955000 ;
      RECT 2.990000  0.295000 3.420000 0.465000 ;
      RECT 3.150000  1.490000 3.420000 1.660000 ;
      RECT 3.150000  1.660000 3.320000 1.785000 ;
      RECT 3.250000  0.465000 3.420000 1.060000 ;
      RECT 3.250000  1.060000 3.485000 1.390000 ;
      RECT 3.250000  1.390000 3.420000 1.490000 ;
      RECT 3.310000  2.125000 3.825000 2.295000 ;
      RECT 3.575000  1.810000 3.825000 2.125000 ;
      RECT 3.590000  0.345000 3.825000 0.675000 ;
      RECT 3.655000  0.675000 3.825000 1.810000 ;
      RECT 3.995000  0.345000 4.185000 2.125000 ;
      RECT 3.995000  2.125000 4.520000 2.295000 ;
      RECT 4.400000  0.255000 4.605000 0.585000 ;
      RECT 4.400000  0.585000 4.570000 1.565000 ;
      RECT 4.400000  1.565000 5.500000 1.735000 ;
      RECT 4.400000  1.735000 4.590000 1.895000 ;
      RECT 4.760000  2.005000 5.105000 2.635000 ;
      RECT 4.800000  0.085000 5.130000 0.545000 ;
      RECT 5.330000  0.295000 6.225000 0.465000 ;
      RECT 5.330000  0.465000 5.500000 1.565000 ;
      RECT 5.330000  1.735000 5.500000 2.155000 ;
      RECT 5.330000  2.155000 6.280000 2.325000 ;
      RECT 5.670000  0.705000 6.290000 1.035000 ;
      RECT 5.670000  1.035000 5.960000 1.985000 ;
      RECT 6.530000  2.125000 6.850000 2.295000 ;
      RECT 6.680000  1.495000 7.290000 1.665000 ;
      RECT 6.680000  1.665000 6.850000 2.125000 ;
      RECT 7.020000  0.085000 7.270000 0.815000 ;
      RECT 7.020000  1.835000 7.190000 2.635000 ;
      RECT 7.120000  0.995000 7.430000 1.325000 ;
      RECT 7.120000  1.325000 7.290000 1.495000 ;
      RECT 7.940000  0.085000 8.190000 0.885000 ;
      RECT 7.940000  1.495000 8.190000 2.635000 ;
      RECT 8.855000  0.085000 9.105000 0.885000 ;
      RECT 8.855000  1.495000 9.105000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.530000  1.785000 1.700000 1.955000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 1.990000  2.125000 2.160000 2.295000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.370000  2.125000 3.540000 2.295000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.290000  2.125000 4.460000 2.295000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.670000  1.785000 5.840000 1.955000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.590000  2.125000 6.760000 2.295000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
    LAYER met1 ;
      RECT 1.470000 1.755000 1.760000 1.800000 ;
      RECT 1.470000 1.800000 5.900000 1.940000 ;
      RECT 1.470000 1.940000 1.760000 1.985000 ;
      RECT 1.930000 2.095000 2.220000 2.140000 ;
      RECT 1.930000 2.140000 3.600000 2.280000 ;
      RECT 1.930000 2.280000 2.220000 2.325000 ;
      RECT 3.310000 2.095000 3.600000 2.140000 ;
      RECT 3.310000 2.280000 3.600000 2.325000 ;
      RECT 4.230000 2.095000 4.520000 2.140000 ;
      RECT 4.230000 2.140000 6.820000 2.280000 ;
      RECT 4.230000 2.280000 4.520000 2.325000 ;
      RECT 5.610000 1.755000 5.900000 1.800000 ;
      RECT 5.610000 1.940000 5.900000 1.985000 ;
      RECT 6.530000 2.095000 6.820000 2.140000 ;
      RECT 6.530000 2.280000 6.820000 2.325000 ;
  END
END sky130_fd_sc_hd__mux4_4
MACRO sky130_fd_sc_hd__nand2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.940000 1.075000 1.275000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.055000 0.430000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 1.485000 0.865000 2.465000 ;
        RECT 0.600000 0.255000 1.295000 0.885000 ;
        RECT 0.600000 0.885000 0.770000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.085000 0.310000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.085000  0.085000 0.395000 0.885000 ;
      RECT 0.085000  1.495000 0.365000 2.635000 ;
      RECT 1.035000  1.495000 1.295000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__nand2_1
MACRO sky130_fd_sc_hd__nand2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 1.075000 1.765000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.845000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.495000 2.215000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 0.655000 2.215000 0.905000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
        RECT 1.935000 0.905000 2.215000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.085000  0.255000 0.425000 0.715000 ;
      RECT 0.085000  0.715000 1.185000 0.885000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.545000 ;
      RECT 0.935000  0.255000 2.105000 0.465000 ;
      RECT 0.935000  0.465000 1.185000 0.715000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.775000  0.465000 2.105000 0.485000 ;
      RECT 1.855000  1.835000 2.110000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__nand2_2
MACRO sky130_fd_sc_hd__nand2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615000 1.075000 4.055000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 1.730000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.495000 3.365000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
        RECT 1.910000 1.075000 2.445000 1.495000 ;
        RECT 2.195000 0.635000 3.365000 0.805000 ;
        RECT 2.195000 0.805000 2.445000 1.075000 ;
        RECT 2.195000 1.665000 2.525000 2.465000 ;
        RECT 3.035000 1.665000 3.365000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.715000 ;
      RECT 0.090000  0.715000 2.025000 0.905000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.545000 ;
      RECT 0.935000  0.255000 1.265000 0.715000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.435000  0.085000 1.605000 0.545000 ;
      RECT 1.775000  0.255000 3.785000 0.465000 ;
      RECT 1.775000  0.465000 2.025000 0.715000 ;
      RECT 1.855000  1.835000 2.025000 2.635000 ;
      RECT 2.695000  1.835000 2.865000 2.635000 ;
      RECT 3.535000  0.465000 3.785000 0.885000 ;
      RECT 3.535000  1.835000 3.785000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__nand2_4
MACRO sky130_fd_sc_hd__nand2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.290000 1.075000 6.305000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.510000 1.075000 3.365000 1.295000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  2.862000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.465000 6.725000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
        RECT 2.195000 1.665000 2.525000 2.465000 ;
        RECT 3.035000 1.665000 3.365000 2.465000 ;
        RECT 3.640000 1.075000 4.120000 1.465000 ;
        RECT 3.875000 0.655000 6.725000 0.905000 ;
        RECT 3.875000 0.905000 4.120000 1.075000 ;
        RECT 3.875000 1.665000 4.205000 2.465000 ;
        RECT 4.715000 1.665000 5.045000 2.465000 ;
        RECT 5.555000 1.665000 5.885000 2.465000 ;
        RECT 6.395000 1.665000 6.725000 2.465000 ;
        RECT 6.475000 0.905000 6.725000 1.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.735000 ;
      RECT 0.090000  0.735000 3.705000 0.905000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.565000 ;
      RECT 0.935000  0.255000 1.265000 0.735000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.435000  0.085000 1.605000 0.565000 ;
      RECT 1.775000  0.255000 2.105000 0.735000 ;
      RECT 1.855000  1.835000 2.025000 2.635000 ;
      RECT 2.275000  0.085000 2.445000 0.565000 ;
      RECT 2.615000  0.255000 2.945000 0.735000 ;
      RECT 2.695000  1.835000 2.865000 2.635000 ;
      RECT 3.115000  0.085000 3.285000 0.565000 ;
      RECT 3.455000  0.255000 7.270000 0.485000 ;
      RECT 3.455000  0.485000 3.705000 0.735000 ;
      RECT 3.535000  1.835000 3.705000 2.635000 ;
      RECT 4.375000  1.835000 4.545000 2.635000 ;
      RECT 5.215000  1.835000 5.385000 2.635000 ;
      RECT 6.055000  1.835000 6.225000 2.635000 ;
      RECT 6.895000  0.485000 7.270000 0.905000 ;
      RECT 6.915000  1.495000 7.270000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__nand2_8
MACRO sky130_fd_sc_hd__nand2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.440000 1.315000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 1.075000 1.085000 1.315000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 1.835000 2.170000 2.005000 ;
        RECT 1.000000 2.005000 1.330000 2.465000 ;
        RECT 1.420000 0.255000 2.170000 0.545000 ;
        RECT 1.800000 0.545000 2.170000 1.835000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.090000  0.525000 0.360000 0.735000 ;
      RECT 0.090000  0.735000 1.425000 0.905000 ;
      RECT 0.090000  1.495000 1.425000 1.665000 ;
      RECT 0.090000  1.665000 0.370000 1.825000 ;
      RECT 0.580000  0.085000 0.910000 0.545000 ;
      RECT 0.580000  1.835000 0.830000 2.635000 ;
      RECT 1.255000  0.905000 1.425000 1.075000 ;
      RECT 1.255000  1.075000 1.630000 1.325000 ;
      RECT 1.255000  1.325000 1.425000 1.495000 ;
      RECT 1.500000  2.175000 1.715000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__nand2b_1
MACRO sky130_fd_sc_hd__nand2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 0.995000 0.800000 1.325000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 1.075000 3.135000 1.275000 ;
        RECT 1.990000 1.275000 2.180000 1.655000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.775500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 1.835000 2.635000 2.005000 ;
        RECT 1.035000 2.005000 1.365000 2.465000 ;
        RECT 1.525000 0.635000 1.855000 0.805000 ;
        RECT 1.530000 0.805000 1.855000 0.905000 ;
        RECT 1.530000 0.905000 1.810000 1.835000 ;
        RECT 2.280000 2.005000 2.635000 2.465000 ;
        RECT 2.360000 1.495000 2.635000 1.835000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.110000  0.510000 0.345000 0.840000 ;
      RECT 0.110000  0.840000 0.280000 1.495000 ;
      RECT 0.110000  1.495000 1.360000 1.665000 ;
      RECT 0.110000  1.665000 0.410000 1.860000 ;
      RECT 0.515000  0.085000 0.845000 0.825000 ;
      RECT 0.580000  1.835000 0.835000 2.635000 ;
      RECT 1.030000  1.075000 1.360000 1.495000 ;
      RECT 1.080000  0.255000 2.275000 0.465000 ;
      RECT 1.080000  0.465000 1.355000 0.905000 ;
      RECT 1.535000  2.175000 2.110000 2.635000 ;
      RECT 2.025000  0.465000 2.275000 0.695000 ;
      RECT 2.025000  0.695000 3.135000 0.905000 ;
      RECT 2.445000  0.085000 2.615000 0.525000 ;
      RECT 2.785000  0.255000 3.135000 0.695000 ;
      RECT 2.805000  1.495000 3.135000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__nand2b_2
MACRO sky130_fd_sc_hd__nand2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.155000 1.075000 4.940000 1.275000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.635000 2.640000 0.905000 ;
        RECT 1.455000 1.445000 4.320000 1.665000 ;
        RECT 1.455000 1.665000 1.785000 2.465000 ;
        RECT 2.295000 1.665000 2.640000 2.465000 ;
        RECT 2.375000 0.905000 2.640000 1.445000 ;
        RECT 3.150000 1.665000 3.480000 2.465000 ;
        RECT 3.990000 1.665000 4.320000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.715000 ;
      RECT 0.090000  0.715000 0.780000 0.905000 ;
      RECT 0.090000  1.445000 0.780000 1.665000 ;
      RECT 0.090000  1.665000 0.425000 2.465000 ;
      RECT 0.595000  0.085000 0.790000 0.545000 ;
      RECT 0.595000  1.835000 1.285000 2.635000 ;
      RECT 0.610000  0.905000 0.780000 1.075000 ;
      RECT 0.610000  1.075000 2.205000 1.275000 ;
      RECT 0.610000  1.275000 0.780000 1.445000 ;
      RECT 0.970000  1.445000 1.285000 1.835000 ;
      RECT 1.035000  0.255000 3.060000 0.465000 ;
      RECT 1.035000  0.465000 1.285000 0.905000 ;
      RECT 1.955000  1.835000 2.125000 2.635000 ;
      RECT 2.810000  0.465000 3.060000 0.715000 ;
      RECT 2.810000  0.715000 4.850000 0.905000 ;
      RECT 2.810000  1.835000 2.980000 2.635000 ;
      RECT 3.230000  0.085000 3.400000 0.545000 ;
      RECT 3.570000  0.255000 3.900000 0.715000 ;
      RECT 3.650000  1.835000 3.820000 2.635000 ;
      RECT 4.070000  0.085000 4.310000 0.545000 ;
      RECT 4.520000  0.255000 4.850000 0.715000 ;
      RECT 4.520000  1.495000 4.850000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__nand2b_4
MACRO sky130_fd_sc_hd__nand3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445000 0.995000 1.755000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 0.765000 1.240000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 0.745000 0.330000 1.325000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.699000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 1.745000 0.595000 ;
        RECT 0.515000 0.595000 0.695000 1.495000 ;
        RECT 0.515000 1.495000 1.745000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.415000 0.595000 1.745000 0.825000 ;
        RECT 1.415000 1.665000 1.745000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.090000  0.085000 0.345000 0.575000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 1.015000  1.835000 1.245000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__nand3_1
MACRO sky130_fd_sc_hd__nand3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.330000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 1.075000 2.160000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.470000 1.075000 3.595000 1.275000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.985500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.635000 0.845000 1.445000 ;
        RECT 0.515000 1.445000 3.045000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
        RECT 2.715000 1.665000 3.045000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.090000  0.295000 2.105000 0.465000 ;
      RECT 0.090000  0.465000 0.345000 0.785000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.355000  0.635000 3.045000 0.905000 ;
      RECT 1.855000  1.835000 2.545000 2.635000 ;
      RECT 2.295000  0.085000 2.625000 0.465000 ;
      RECT 3.215000  0.085000 3.595000 0.885000 ;
      RECT 3.215000  1.445000 3.595000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__nand3_2
MACRO sky130_fd_sc_hd__nand3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.850000 1.075000 5.565000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 1.075000 3.540000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 1.700000 1.275000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.971000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.445000 6.355000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
        RECT 2.195000 1.665000 2.525000 2.465000 ;
        RECT 3.035000 1.665000 3.365000 2.465000 ;
        RECT 4.395000 0.655000 6.355000 0.905000 ;
        RECT 4.395000 1.665000 4.725000 2.465000 ;
        RECT 5.235000 1.665000 5.565000 2.465000 ;
        RECT 6.125000 0.905000 6.355000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.735000 ;
      RECT 0.090000  0.735000 3.785000 0.905000 ;
      RECT 0.090000  1.445000 0.345000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.565000 ;
      RECT 0.935000  0.255000 1.265000 0.735000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.435000  0.085000 1.605000 0.565000 ;
      RECT 1.775000  0.655000 2.105000 0.735000 ;
      RECT 1.855000  1.835000 2.025000 2.635000 ;
      RECT 2.195000  0.255000 6.000000 0.485000 ;
      RECT 2.615000  0.655000 2.945000 0.735000 ;
      RECT 2.695000  1.835000 2.865000 2.635000 ;
      RECT 3.455000  0.655000 3.785000 0.735000 ;
      RECT 3.535000  1.835000 4.225000 2.635000 ;
      RECT 4.895000  1.835000 5.065000 2.635000 ;
      RECT 5.735000  1.835000 6.000000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__nand3_4
MACRO sky130_fd_sc_hd__nand3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.325000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.425000 0.995000 1.755000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 0.995000 1.235000 1.325000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.732000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.130000 1.495000 2.675000 1.665000 ;
        RECT 1.130000 1.665000 1.460000 2.465000 ;
        RECT 2.085000 0.255000 2.675000 0.485000 ;
        RECT 2.085000 1.665000 2.675000 2.465000 ;
        RECT 2.385000 0.485000 2.675000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.445000 0.510000 0.655000 ;
      RECT 0.085000  0.655000 2.215000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.595000 ;
      RECT 0.085000  1.595000 0.510000 1.925000 ;
      RECT 0.710000  0.085000 1.040000 0.485000 ;
      RECT 0.710000  1.495000 0.960000 2.635000 ;
      RECT 1.630000  1.835000 1.915000 2.635000 ;
      RECT 2.045000  0.825000 2.215000 1.325000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__nand3b_1
MACRO sky130_fd_sc_hd__nand3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.075000 0.780000 1.275000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.950000 1.075000 3.140000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 1.075000 1.740000 1.275000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.985500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 1.785000 4.050000 1.955000 ;
        RECT 1.060000 1.955000 2.230000 2.005000 ;
        RECT 1.060000 2.005000 1.390000 2.465000 ;
        RECT 1.900000 2.005000 2.230000 2.465000 ;
        RECT 3.260000 0.635000 4.050000 0.905000 ;
        RECT 3.260000 1.955000 4.050000 2.005000 ;
        RECT 3.260000 2.005000 3.510000 2.465000 ;
        RECT 3.850000 0.905000 4.050000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.255000 0.410000 0.655000 ;
      RECT 0.090000  0.655000 0.260000 1.445000 ;
      RECT 0.090000  1.445000 3.650000 1.615000 ;
      RECT 0.090000  1.615000 0.260000 2.065000 ;
      RECT 0.090000  2.065000 0.410000 2.465000 ;
      RECT 0.580000  0.085000 0.890000 0.905000 ;
      RECT 0.580000  1.835000 0.890000 2.635000 ;
      RECT 1.060000  0.255000 1.390000 0.715000 ;
      RECT 1.060000  0.715000 2.750000 0.905000 ;
      RECT 1.560000  0.085000 1.810000 0.545000 ;
      RECT 1.560000  2.175000 1.730000 2.635000 ;
      RECT 2.000000  0.255000 4.050000 0.465000 ;
      RECT 2.000000  0.635000 2.750000 0.715000 ;
      RECT 2.400000  2.175000 2.650000 2.635000 ;
      RECT 2.840000  2.175000 3.090000 2.635000 ;
      RECT 2.920000  0.465000 3.090000 0.905000 ;
      RECT 3.320000  1.075000 3.650000 1.445000 ;
      RECT 3.760000  2.175000 4.050000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__nand3b_2
MACRO sky130_fd_sc_hd__nand3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.075000 0.780000 1.275000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.270000 1.075000 4.480000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.790000 1.075000 6.500000 1.275000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.971000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.635000 2.965000 0.905000 ;
        RECT 1.455000 1.445000 6.505000 1.665000 ;
        RECT 1.455000 1.665000 1.785000 2.465000 ;
        RECT 2.295000 1.665000 3.465000 2.005000 ;
        RECT 2.295000 2.005000 2.625000 2.465000 ;
        RECT 2.795000 0.905000 2.965000 1.075000 ;
        RECT 2.795000 1.075000 3.100000 1.445000 ;
        RECT 3.135000 2.005000 3.465000 2.465000 ;
        RECT 3.975000 1.665000 4.305000 2.465000 ;
        RECT 5.335000 1.665000 5.665000 2.465000 ;
        RECT 6.175000 1.665000 6.505000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.085000  0.255000 0.425000 0.715000 ;
      RECT 0.085000  0.715000 1.285000 0.905000 ;
      RECT 0.085000  0.905000 0.260000 1.445000 ;
      RECT 0.085000  1.445000 0.425000 2.465000 ;
      RECT 0.595000  0.085000 0.845000 0.545000 ;
      RECT 0.595000  1.445000 1.285000 2.635000 ;
      RECT 1.005000  0.905000 1.285000 1.075000 ;
      RECT 1.005000  1.075000 2.625000 1.275000 ;
      RECT 1.035000  0.255000 4.725000 0.465000 ;
      RECT 1.955000  1.835000 2.125000 2.635000 ;
      RECT 2.795000  2.175000 2.965000 2.635000 ;
      RECT 3.135000  0.635000 4.725000 0.715000 ;
      RECT 3.135000  0.715000 6.505000 0.905000 ;
      RECT 3.635000  1.835000 3.805000 2.635000 ;
      RECT 4.475000  1.835000 5.165000 2.635000 ;
      RECT 4.915000  0.085000 5.165000 0.545000 ;
      RECT 5.335000  0.255000 5.665000 0.715000 ;
      RECT 5.835000  0.085000 6.005000 0.545000 ;
      RECT 5.835000  1.835000 6.005000 2.635000 ;
      RECT 6.175000  0.255000 6.505000 0.715000 ;
      RECT 6.675000  0.085000 7.005000 0.905000 ;
      RECT 6.675000  1.445000 7.005000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__nand3b_4
MACRO sky130_fd_sc_hd__nand4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 0.995000 2.215000 1.665000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 0.300000 1.350000 0.825000 ;
        RECT 1.145000 0.825000 1.350000 0.995000 ;
        RECT 1.145000 0.995000 1.455000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.300000 0.810000 0.995000 ;
        RECT 0.595000 0.995000 0.975000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 0.995000 0.395000 1.325000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.795000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.495000 1.795000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.385000 1.665000 1.715000 2.465000 ;
        RECT 1.520000 0.255000 2.215000 0.825000 ;
        RECT 1.625000 0.825000 1.795000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 0.090000  0.085000 0.425000 0.825000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.915000  1.835000 2.195000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__nand4_1
MACRO sky130_fd_sc_hd__nand4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165000 1.075000 4.495000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.235000 1.075000 3.080000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 1.075000 1.700000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.845000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.255500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.445000 3.925000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
        RECT 2.355000 1.665000 2.685000 2.465000 ;
        RECT 3.370000 1.055000 3.925000 1.445000 ;
        RECT 3.595000 0.635000 3.925000 1.055000 ;
        RECT 3.595000 1.665000 3.925000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.735000 ;
      RECT 0.090000  0.735000 1.185000 0.905000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.545000 ;
      RECT 0.935000  0.255000 2.125000 0.465000 ;
      RECT 0.935000  0.465000 1.185000 0.735000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.355000  0.635000 3.085000 0.905000 ;
      RECT 1.855000  1.835000 2.185000 2.635000 ;
      RECT 2.315000  0.255000 4.425000 0.465000 ;
      RECT 2.995000  1.835000 3.325000 2.635000 ;
      RECT 3.255000  0.465000 3.425000 0.885000 ;
      RECT 4.095000  0.465000 4.425000 0.905000 ;
      RECT 4.095000  1.445000 4.425000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__nand4_2
MACRO sky130_fd_sc_hd__nand4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.465000 1.075000 7.710000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.850000 1.075000 5.565000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 1.075000 3.540000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 1.700000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.511000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.445000 7.305000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
        RECT 2.195000 1.665000 2.525000 2.465000 ;
        RECT 3.035000 1.665000 3.365000 2.465000 ;
        RECT 4.395000 1.665000 4.725000 2.465000 ;
        RECT 5.235000 1.665000 5.565000 2.465000 ;
        RECT 6.110000 0.655000 7.305000 0.905000 ;
        RECT 6.110000 0.905000 6.290000 1.445000 ;
        RECT 6.135000 1.665000 6.465000 2.465000 ;
        RECT 6.975000 1.665000 7.305000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.090000  0.255000 0.345000 0.655000 ;
      RECT 0.090000  0.655000 2.025000 0.905000 ;
      RECT 0.090000  1.445000 0.345000 2.635000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 1.015000  0.255000 1.185000 0.655000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.355000  0.085000 1.685000 0.485000 ;
      RECT 1.855000  0.255000 3.785000 0.485000 ;
      RECT 1.855000  0.485000 2.025000 0.655000 ;
      RECT 1.855000  1.835000 2.025000 2.635000 ;
      RECT 2.195000  0.655000 5.565000 0.905000 ;
      RECT 2.695000  1.835000 2.865000 2.635000 ;
      RECT 3.535000  1.835000 4.225000 2.635000 ;
      RECT 3.975000  0.255000 7.730000 0.485000 ;
      RECT 4.895000  1.835000 5.065000 2.635000 ;
      RECT 5.770000  0.485000 5.940000 0.905000 ;
      RECT 5.770000  1.835000 5.940000 2.635000 ;
      RECT 6.635000  1.835000 6.805000 2.635000 ;
      RECT 7.475000  0.485000 7.730000 0.905000 ;
      RECT 7.475000  1.445000 7.735000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__nand4_4
MACRO sky130_fd_sc_hd__nand4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.325000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925000 0.765000 2.185000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 0.765000 1.755000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 0.995000 1.235000 1.325000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.887500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.130000 1.495000 3.135000 1.665000 ;
        RECT 1.130000 1.665000 1.460000 2.465000 ;
        RECT 2.085000 1.665000 2.415000 2.465000 ;
        RECT 2.695000 0.255000 3.135000 0.825000 ;
        RECT 2.925000 0.825000 3.135000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.445000 0.475000 0.655000 ;
      RECT 0.085000  0.655000 1.335000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.595000 ;
      RECT 0.085000  1.595000 0.510000 1.925000 ;
      RECT 0.655000  0.085000 0.985000 0.485000 ;
      RECT 0.710000  1.495000 0.960000 2.635000 ;
      RECT 1.155000  0.425000 2.525000 0.595000 ;
      RECT 1.155000  0.595000 1.335000 0.655000 ;
      RECT 1.630000  1.835000 1.915000 2.635000 ;
      RECT 2.355000  0.595000 2.525000 0.995000 ;
      RECT 2.355000  0.995000 2.755000 1.325000 ;
      RECT 2.705000  1.835000 2.920000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__nand4b_1
MACRO sky130_fd_sc_hd__nand4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.330000 1.615000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.010000 1.075000 3.100000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.360000 1.075000 4.450000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.620000 1.075000 5.430000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.255500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.635000 1.785000 0.825000 ;
        RECT 1.455000 1.445000 4.865000 1.665000 ;
        RECT 1.455000 1.665000 1.785000 2.465000 ;
        RECT 1.550000 0.825000 1.785000 1.445000 ;
        RECT 2.295000 1.665000 2.625000 2.465000 ;
        RECT 3.605000 1.665000 3.935000 2.465000 ;
        RECT 4.535000 1.665000 4.865000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.090000  0.255000 0.345000 0.635000 ;
      RECT 0.090000  0.635000 0.670000 0.805000 ;
      RECT 0.090000  1.915000 0.670000 2.085000 ;
      RECT 0.090000  2.085000 0.345000 2.465000 ;
      RECT 0.500000  0.805000 0.670000 1.075000 ;
      RECT 0.500000  1.075000 1.380000 1.245000 ;
      RECT 0.500000  1.245000 0.670000 1.915000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.255000 1.285000 2.635000 ;
      RECT 1.035000  0.255000 2.125000 0.465000 ;
      RECT 1.035000  0.465000 1.285000 0.905000 ;
      RECT 1.035000  1.445000 1.285000 2.255000 ;
      RECT 1.955000  0.465000 2.125000 0.635000 ;
      RECT 1.955000  0.635000 3.045000 0.905000 ;
      RECT 1.955000  1.835000 2.125000 2.635000 ;
      RECT 2.295000  0.255000 3.985000 0.465000 ;
      RECT 2.795000  1.835000 3.435000 2.635000 ;
      RECT 3.235000  0.635000 4.455000 0.715000 ;
      RECT 3.235000  0.715000 5.340000 0.905000 ;
      RECT 4.105000  1.835000 4.365000 2.635000 ;
      RECT 4.155000  0.255000 4.415000 0.615000 ;
      RECT 4.155000  0.615000 4.455000 0.635000 ;
      RECT 4.665000  0.085000 4.835000 0.545000 ;
      RECT 5.005000  0.255000 5.340000 0.715000 ;
      RECT 5.035000  1.495000 5.430000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__nand4b_2
MACRO sky130_fd_sc_hd__nand4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.930000 1.075000 4.590000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.790000 1.075000 6.510000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.015000 1.075000 8.655000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.511000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.635000 2.640000 0.905000 ;
        RECT 1.455000 1.445000 8.185000 1.665000 ;
        RECT 1.455000 1.665000 1.785000 2.465000 ;
        RECT 2.295000 1.665000 2.625000 2.465000 ;
        RECT 2.375000 0.905000 2.640000 1.445000 ;
        RECT 3.135000 1.665000 3.465000 2.465000 ;
        RECT 3.975000 1.665000 4.305000 2.465000 ;
        RECT 5.335000 1.665000 5.665000 2.465000 ;
        RECT 6.175000 1.665000 6.505000 2.465000 ;
        RECT 7.015000 1.665000 7.345000 2.465000 ;
        RECT 7.855000 1.665000 8.185000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.930000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.735000 ;
      RECT 0.090000  0.735000 0.805000 0.905000 ;
      RECT 0.090000  1.495000 0.805000 1.665000 ;
      RECT 0.090000  1.665000 0.425000 2.465000 ;
      RECT 0.595000  0.085000 0.845000 0.545000 ;
      RECT 0.595000  1.835000 1.285000 2.635000 ;
      RECT 0.610000  0.905000 0.805000 1.075000 ;
      RECT 0.610000  1.075000 2.205000 1.275000 ;
      RECT 0.610000  1.275000 0.805000 1.495000 ;
      RECT 0.995000  1.495000 1.285000 1.835000 ;
      RECT 1.035000  0.255000 4.725000 0.465000 ;
      RECT 1.035000  0.465000 1.285000 0.905000 ;
      RECT 1.955000  1.835000 2.125000 2.635000 ;
      RECT 2.795000  1.835000 2.965000 2.635000 ;
      RECT 3.135000  0.635000 6.505000 0.905000 ;
      RECT 3.635000  1.835000 3.805000 2.635000 ;
      RECT 4.475000  1.835000 5.165000 2.635000 ;
      RECT 4.915000  0.255000 6.925000 0.465000 ;
      RECT 5.835000  1.835000 6.005000 2.635000 ;
      RECT 6.675000  0.465000 6.925000 0.735000 ;
      RECT 6.675000  0.735000 8.610000 0.905000 ;
      RECT 6.675000  1.835000 6.845000 2.635000 ;
      RECT 7.095000  0.085000 7.265000 0.545000 ;
      RECT 7.435000  0.255000 7.765000 0.735000 ;
      RECT 7.515000  1.835000 7.685000 2.635000 ;
      RECT 7.935000  0.085000 8.105000 0.545000 ;
      RECT 8.275000  0.255000 8.610000 0.735000 ;
      RECT 8.355000  1.445000 8.610000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
  END
END sky130_fd_sc_hd__nand4b_4
MACRO sky130_fd_sc_hd__nand4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.390000 0.725000 3.640000 1.615000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.075000 0.780000 1.655000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 0.735000 1.720000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.970000 1.075000 1.320000 1.325000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.909000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.120000 1.495000 2.670000 1.665000 ;
        RECT 1.120000 1.665000 1.450000 2.465000 ;
        RECT 2.140000 1.665000 2.470000 2.465000 ;
        RECT 2.420000 0.255000 2.930000 0.825000 ;
        RECT 2.420000 0.825000 2.670000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.485000 0.425000 0.715000 ;
      RECT 0.085000  0.715000 1.270000 0.905000 ;
      RECT 0.085000  0.905000 0.260000 2.065000 ;
      RECT 0.085000  2.065000 0.425000 2.465000 ;
      RECT 0.595000  0.085000 0.900000 0.545000 ;
      RECT 0.595000  1.835000 0.925000 2.635000 ;
      RECT 1.080000  0.365000 2.250000 0.555000 ;
      RECT 1.080000  0.555000 1.270000 0.715000 ;
      RECT 1.640000  1.835000 1.970000 2.635000 ;
      RECT 1.970000  0.555000 2.250000 1.325000 ;
      RECT 2.680000  2.175000 3.450000 2.635000 ;
      RECT 2.840000  0.995000 3.090000 1.835000 ;
      RECT 2.840000  1.835000 4.055000 2.005000 ;
      RECT 3.100000  0.085000 3.450000 0.545000 ;
      RECT 3.620000  0.255000 4.055000 0.545000 ;
      RECT 3.635000  2.005000 4.055000 2.465000 ;
      RECT 3.810000  0.545000 4.055000 1.835000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__nand4bb_1
MACRO sky130_fd_sc_hd__nand4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.170000 0.890000 1.340000 ;
        RECT 0.610000 1.070000 0.890000 1.170000 ;
        RECT 0.610000 1.340000 0.890000 1.615000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.070000 0.330000 1.615000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.720000 1.075000 4.615000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.945000 1.075000 5.875000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.255500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.085000 0.655000 2.415000 1.445000 ;
        RECT 2.085000 1.445000 5.455000 1.665000 ;
        RECT 2.085000 1.665000 2.335000 2.465000 ;
        RECT 2.925000 1.665000 3.255000 2.465000 ;
        RECT 3.245000 1.075000 3.550000 1.445000 ;
        RECT 4.285000 1.665000 4.615000 2.465000 ;
        RECT 5.125000 1.665000 5.455000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.730000 ;
      RECT 0.085000  0.730000 1.230000 0.900000 ;
      RECT 0.085000  1.785000 1.230000 1.980000 ;
      RECT 0.085000  1.980000 0.370000 2.440000 ;
      RECT 0.515000  0.085000 0.765000 0.545000 ;
      RECT 0.540000  2.195000 0.765000 2.635000 ;
      RECT 0.935000  0.255000 1.575000 0.560000 ;
      RECT 0.935000  2.150000 1.575000 2.465000 ;
      RECT 1.060000  0.900000 1.230000 1.785000 ;
      RECT 1.400000  0.560000 1.575000 0.715000 ;
      RECT 1.400000  0.715000 1.580000 1.410000 ;
      RECT 1.400000  1.410000 1.575000 2.150000 ;
      RECT 1.745000  0.255000 3.675000 0.485000 ;
      RECT 1.745000  0.485000 1.915000 0.585000 ;
      RECT 1.745000  1.495000 1.915000 2.635000 ;
      RECT 2.505000  1.835000 2.755000 2.635000 ;
      RECT 2.745000  1.075000 3.075000 1.275000 ;
      RECT 2.925000  0.655000 4.615000 0.905000 ;
      RECT 3.425000  1.835000 4.115000 2.635000 ;
      RECT 3.865000  0.255000 5.035000 0.485000 ;
      RECT 4.785000  0.485000 5.035000 0.735000 ;
      RECT 4.785000  0.735000 5.895000 0.905000 ;
      RECT 4.785000  1.835000 4.955000 2.635000 ;
      RECT 5.205000  0.085000 5.375000 0.565000 ;
      RECT 5.545000  0.255000 5.895000 0.735000 ;
      RECT 5.625000  1.445000 5.895000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.060000  1.105000 1.230000 1.275000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  1.105000 3.075000 1.275000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 1.000000 1.075000 3.135000 1.305000 ;
  END
END sky130_fd_sc_hd__nand4bb_2
MACRO sky130_fd_sc_hd__nand4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.995000 0.330000 1.615000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.590000 0.995000 0.975000 1.615000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.120000 1.075000 7.910000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.420000 1.075000 10.015000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.511000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.540000 0.655000 3.990000 0.905000 ;
        RECT 2.540000 1.445000 9.590000 1.665000 ;
        RECT 2.540000 1.665000 2.790000 2.465000 ;
        RECT 3.380000 1.665000 3.710000 2.465000 ;
        RECT 3.700000 0.905000 3.990000 1.445000 ;
        RECT 4.220000 1.665000 4.550000 2.465000 ;
        RECT 5.060000 1.665000 5.390000 2.465000 ;
        RECT 6.740000 1.665000 7.070000 2.465000 ;
        RECT 7.580000 1.665000 7.910000 2.465000 ;
        RECT 8.420000 1.665000 8.750000 2.465000 ;
        RECT 9.260000 1.665000 9.590000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.085000  0.255000  0.345000 0.635000 ;
      RECT 0.085000  0.635000  1.455000 0.805000 ;
      RECT 0.085000  1.785000  1.455000 1.980000 ;
      RECT 0.085000  1.980000  0.370000 2.440000 ;
      RECT 0.515000  0.085000  0.845000 0.465000 ;
      RECT 0.540000  2.195000  0.765000 2.635000 ;
      RECT 0.935000  2.150000  1.795000 2.465000 ;
      RECT 1.015000  0.255000  1.795000 0.465000 ;
      RECT 1.145000  0.805000  1.455000 1.785000 ;
      RECT 1.625000  0.465000  1.795000 1.075000 ;
      RECT 1.625000  1.075000  2.210000 1.305000 ;
      RECT 1.625000  1.305000  1.795000 2.150000 ;
      RECT 2.200000  0.255000  5.810000 0.485000 ;
      RECT 2.200000  0.485000  2.370000 0.905000 ;
      RECT 2.200000  1.495000  2.370000 2.635000 ;
      RECT 2.540000  1.075000  3.285000 1.245000 ;
      RECT 2.960000  1.835000  3.210000 2.635000 ;
      RECT 3.880000  1.835000  4.050000 2.635000 ;
      RECT 4.160000  1.075000  5.390000 1.275000 ;
      RECT 4.220000  0.655000  5.390000 0.735000 ;
      RECT 4.220000  0.735000  6.150000 0.905000 ;
      RECT 4.720000  1.835000  4.890000 2.635000 ;
      RECT 5.610000  1.835000  6.540000 2.635000 ;
      RECT 5.980000  0.255000  7.910000 0.485000 ;
      RECT 5.980000  0.485000  6.150000 0.735000 ;
      RECT 6.320000  0.655000 10.035000 0.905000 ;
      RECT 7.240000  1.835000  7.410000 2.635000 ;
      RECT 8.080000  1.835000  8.250000 2.635000 ;
      RECT 8.420000  0.085000  8.750000 0.485000 ;
      RECT 8.920000  1.835000  9.090000 2.635000 ;
      RECT 9.260000  0.085000  9.590000 0.485000 ;
      RECT 9.760000  1.445000 10.035000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.980000  1.105000 2.150000 1.275000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.280000  1.105000 4.450000 1.275000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
    LAYER met1 ;
      RECT 1.920000 1.075000 2.210000 1.120000 ;
      RECT 1.920000 1.120000 4.510000 1.260000 ;
      RECT 1.920000 1.260000 2.210000 1.305000 ;
      RECT 4.220000 1.075000 4.510000 1.120000 ;
      RECT 4.220000 1.260000 4.510000 1.305000 ;
  END
END sky130_fd_sc_hd__nand4bb_4
MACRO sky130_fd_sc_hd__nor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 1.075000 1.295000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.435000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.495000 0.775000 1.665000 ;
        RECT 0.095000 1.665000 0.425000 2.450000 ;
        RECT 0.515000 0.255000 0.845000 0.895000 ;
        RECT 0.605000 0.895000 0.775000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.105000  0.085000 0.345000 0.895000 ;
      RECT 0.955000  1.495000 1.285000 2.635000 ;
      RECT 1.015000  0.085000 1.285000 0.895000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__nor2_1
MACRO sky130_fd_sc_hd__nor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.810000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.980000 1.075000 1.750000 1.275000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 1.705000 0.735000 ;
        RECT 0.535000 0.735000 2.135000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 1.375000 1.445000 2.135000 1.665000 ;
        RECT 1.375000 1.665000 1.705000 2.125000 ;
        RECT 1.920000 0.905000 2.135000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 1.205000 1.665000 ;
      RECT 0.090000  1.665000 0.365000 2.465000 ;
      RECT 0.535000  1.835000 0.865000 2.635000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.035000  1.665000 1.205000 2.295000 ;
      RECT 1.035000  2.295000 2.175000 2.465000 ;
      RECT 1.875000  0.085000 2.165000 0.555000 ;
      RECT 1.875000  1.835000 2.175000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__nor2_2
MACRO sky130_fd_sc_hd__nor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 1.075000 1.800000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.120000 1.075000 3.485000 1.275000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 4.055000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.215000 0.255000 2.545000 0.725000 ;
        RECT 2.295000 1.445000 4.055000 1.745000 ;
        RECT 2.295000 1.745000 2.465000 2.125000 ;
        RECT 3.055000 0.255000 3.385000 0.725000 ;
        RECT 3.135000 1.745000 3.305000 2.125000 ;
        RECT 3.655000 0.905000 4.055000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 2.125000 1.665000 ;
      RECT 0.090000  1.665000 0.365000 2.465000 ;
      RECT 0.535000  1.835000 0.865000 2.635000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.035000  1.665000 1.205000 2.465000 ;
      RECT 1.375000  1.835000 1.625000 2.635000 ;
      RECT 1.795000  1.665000 2.125000 2.295000 ;
      RECT 1.795000  2.295000 3.890000 2.465000 ;
      RECT 1.875000  0.085000 2.045000 0.555000 ;
      RECT 2.635000  1.935000 2.965000 2.295000 ;
      RECT 2.715000  0.085000 2.885000 0.555000 ;
      RECT 3.475000  1.915000 3.890000 2.295000 ;
      RECT 3.555000  0.085000 3.840000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__nor2_4
MACRO sky130_fd_sc_hd__nor2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.360000 1.075000 3.530000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.800000 1.075000 6.540000 1.275000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  2.484000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 7.275000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.215000 0.255000 2.545000 0.725000 ;
        RECT 3.055000 0.255000 3.385000 0.725000 ;
        RECT 3.895000 0.255000 4.225000 0.725000 ;
        RECT 3.935000 1.445000 7.275000 1.615000 ;
        RECT 3.935000 1.615000 4.185000 2.125000 ;
        RECT 4.735000 0.255000 5.065000 0.725000 ;
        RECT 4.775000 1.615000 5.025000 2.125000 ;
        RECT 5.575000 0.255000 5.905000 0.725000 ;
        RECT 5.615000 1.615000 5.865000 2.125000 ;
        RECT 6.415000 0.255000 6.745000 0.725000 ;
        RECT 6.455000 1.615000 6.705000 2.125000 ;
        RECT 6.710000 0.905000 7.275000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 3.765000 1.665000 ;
      RECT 0.090000  1.665000 0.405000 2.465000 ;
      RECT 0.575000  1.835000 0.825000 2.635000 ;
      RECT 0.995000  1.665000 1.245000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.415000  1.835000 1.665000 2.635000 ;
      RECT 1.835000  1.665000 2.085000 2.465000 ;
      RECT 1.875000  0.085000 2.045000 0.555000 ;
      RECT 2.255000  1.835000 2.505000 2.635000 ;
      RECT 2.675000  1.665000 2.925000 2.465000 ;
      RECT 2.715000  0.085000 2.885000 0.555000 ;
      RECT 3.095000  1.835000 3.345000 2.635000 ;
      RECT 3.515000  1.665000 3.765000 2.295000 ;
      RECT 3.515000  2.295000 7.125000 2.465000 ;
      RECT 3.555000  0.085000 3.725000 0.555000 ;
      RECT 4.355000  1.785000 4.605000 2.295000 ;
      RECT 4.395000  0.085000 4.565000 0.555000 ;
      RECT 5.195000  1.785000 5.445000 2.295000 ;
      RECT 5.235000  0.085000 5.405000 0.555000 ;
      RECT 6.035000  1.785000 6.285000 2.295000 ;
      RECT 6.075000  0.085000 6.245000 0.555000 ;
      RECT 6.875000  1.785000 7.125000 2.295000 ;
      RECT 6.915000  0.085000 7.205000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__nor2_8
MACRO sky130_fd_sc_hd__nor2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.960000 1.065000 1.325000 1.325000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.725000 0.325000 1.325000 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.235000 0.255000 1.565000 0.725000 ;
        RECT 1.235000 0.725000 2.215000 0.895000 ;
        RECT 1.655000 1.850000 2.215000 2.465000 ;
        RECT 2.035000 0.895000 2.215000 1.850000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.330000  0.370000 0.675000 0.545000 ;
      RECT 0.415000  1.510000 1.705000 1.680000 ;
      RECT 0.415000  1.680000 0.675000 1.905000 ;
      RECT 0.495000  0.545000 0.675000 1.510000 ;
      RECT 0.855000  0.085000 1.065000 0.895000 ;
      RECT 0.875000  1.855000 1.205000 2.635000 ;
      RECT 1.535000  1.075000 1.865000 1.245000 ;
      RECT 1.535000  1.245000 1.705000 1.510000 ;
      RECT 1.735000  0.085000 2.120000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__nor2b_1
MACRO sky130_fd_sc_hd__nor2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.480000 1.065000 0.920000 1.275000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.600000 1.065000 3.125000 1.275000 ;
        RECT 2.910000 1.275000 3.125000 1.965000 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 1.705000 0.895000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 1.415000 0.895000 1.665000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.085000 0.365000 0.895000 ;
      RECT 0.085000  1.445000 1.245000 1.655000 ;
      RECT 0.085000  1.655000 0.405000 2.465000 ;
      RECT 0.575000  1.825000 0.825000 2.635000 ;
      RECT 0.995000  1.655000 1.245000 2.295000 ;
      RECT 0.995000  2.295000 2.125000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.835000  1.445000 2.090000 1.890000 ;
      RECT 1.835000  1.890000 2.125000 2.295000 ;
      RECT 1.875000  0.085000 2.045000 0.895000 ;
      RECT 1.875000  1.075000 2.430000 1.245000 ;
      RECT 2.215000  0.725000 2.565000 0.895000 ;
      RECT 2.215000  0.895000 2.430000 1.075000 ;
      RECT 2.260000  1.245000 2.430000 1.445000 ;
      RECT 2.260000  1.445000 2.565000 1.615000 ;
      RECT 2.395000  0.445000 2.565000 0.725000 ;
      RECT 2.395000  1.615000 2.565000 2.460000 ;
      RECT 2.775000  0.085000 3.030000 0.845000 ;
      RECT 2.775000  2.145000 3.025000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__nor2b_2
MACRO sky130_fd_sc_hd__nor2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.360000 1.075000 1.800000 1.275000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.075000 4.975000 1.320000 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 3.385000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.215000 0.255000 2.545000 0.725000 ;
        RECT 2.295000 0.905000 2.625000 1.445000 ;
        RECT 2.295000 1.445000 3.305000 1.745000 ;
        RECT 2.295000 1.745000 2.465000 2.125000 ;
        RECT 3.055000 0.255000 3.385000 0.725000 ;
        RECT 3.135000 1.745000 3.305000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.085000 0.365000 0.905000 ;
      RECT 0.085000  1.455000 2.125000 1.665000 ;
      RECT 0.085000  1.665000 0.365000 2.465000 ;
      RECT 0.535000  1.835000 0.865000 2.635000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.035000  1.665000 1.205000 2.465000 ;
      RECT 1.375000  1.835000 1.625000 2.635000 ;
      RECT 1.795000  1.665000 2.125000 2.295000 ;
      RECT 1.795000  2.295000 3.855000 2.465000 ;
      RECT 1.875000  0.085000 2.045000 0.555000 ;
      RECT 2.635000  1.935000 2.965000 2.295000 ;
      RECT 2.715000  0.085000 2.885000 0.555000 ;
      RECT 2.795000  1.075000 4.275000 1.275000 ;
      RECT 3.475000  1.575000 3.855000 2.295000 ;
      RECT 3.555000  0.085000 3.845000 0.905000 ;
      RECT 4.025000  0.255000 4.355000 0.815000 ;
      RECT 4.025000  0.815000 4.275000 1.075000 ;
      RECT 4.025000  1.275000 4.275000 1.575000 ;
      RECT 4.025000  1.575000 4.355000 2.465000 ;
      RECT 4.525000  0.085000 4.815000 0.905000 ;
      RECT 4.525000  1.495000 4.930000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__nor2b_4
MACRO sky130_fd_sc_hd__nor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 0.655000 1.755000 1.665000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.995000 0.975000 1.325000 ;
        RECT 0.595000 1.325000 0.830000 2.005000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.425000 1.325000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.604500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.385000 0.345000 0.655000 ;
        RECT 0.090000 0.655000 1.315000 0.825000 ;
        RECT 0.090000 1.495000 0.425000 2.280000 ;
        RECT 0.090000 2.280000 1.170000 2.450000 ;
        RECT 1.000000 1.495000 1.315000 1.665000 ;
        RECT 1.000000 1.665000 1.170000 2.280000 ;
        RECT 1.015000 0.385000 1.185000 0.655000 ;
        RECT 1.145000 0.825000 1.315000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 1.355000  0.085000 1.685000 0.485000 ;
      RECT 1.435000  1.835000 1.750000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__nor3_1
MACRO sky130_fd_sc_hd__nor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 1.075000 0.965000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135000 1.075000 2.185000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 1.075000 2.965000 1.285000 ;
        RECT 2.375000 1.285000 2.640000 1.625000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.796500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 3.595000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.755000 0.255000 3.085000 0.725000 ;
        RECT 2.835000 1.455000 3.595000 1.625000 ;
        RECT 2.835000 1.625000 3.045000 2.125000 ;
        RECT 3.135000 0.905000 3.595000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.150000  1.455000 2.085000 1.625000 ;
      RECT 0.150000  1.625000 0.405000 2.465000 ;
      RECT 0.575000  1.795000 0.825000 2.635000 ;
      RECT 0.995000  1.625000 1.245000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.415000  1.795000 1.665000 2.295000 ;
      RECT 1.415000  2.295000 3.465000 2.465000 ;
      RECT 1.835000  1.625000 2.085000 2.125000 ;
      RECT 1.875000  0.085000 2.585000 0.555000 ;
      RECT 2.415000  1.795000 2.625000 2.295000 ;
      RECT 3.215000  1.795000 3.465000 2.295000 ;
      RECT 3.255000  0.085000 3.545000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__nor3_2
MACRO sky130_fd_sc_hd__nor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.825000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095000 1.075000 3.685000 1.285000 ;
        RECT 3.515000 1.285000 3.685000 1.445000 ;
        RECT 3.515000 1.445000 5.165000 1.615000 ;
        RECT 4.995000 1.075000 5.415000 1.285000 ;
        RECT 4.995000 1.285000 5.165000 1.445000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.855000 1.075000 4.765000 1.275000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.593000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 5.895000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.215000 0.255000 2.545000 0.725000 ;
        RECT 3.055000 0.255000 3.385000 0.725000 ;
        RECT 3.515000 1.785000 5.895000 1.955000 ;
        RECT 3.515000 1.955000 4.605000 1.965000 ;
        RECT 3.515000 1.965000 3.765000 2.125000 ;
        RECT 3.895000 0.255000 4.225000 0.725000 ;
        RECT 4.355000 1.965000 4.605000 2.125000 ;
        RECT 4.735000 0.255000 5.065000 0.725000 ;
        RECT 5.605000 0.255000 5.895000 0.725000 ;
        RECT 5.605000 0.905000 5.895000 1.785000 ;
        RECT 5.615000 1.955000 5.895000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.150000  1.455000 2.085000 1.625000 ;
      RECT 0.150000  1.625000 0.405000 2.465000 ;
      RECT 0.575000  1.795000 0.825000 2.635000 ;
      RECT 0.995000  1.625000 1.245000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.415000  1.795000 1.665000 2.635000 ;
      RECT 1.835000  1.625000 2.085000 2.085000 ;
      RECT 1.835000  2.085000 2.925000 2.465000 ;
      RECT 1.875000  0.085000 2.045000 0.555000 ;
      RECT 2.255000  1.455000 3.345000 1.625000 ;
      RECT 2.255000  1.625000 2.505000 1.915000 ;
      RECT 2.675000  1.795000 2.925000 2.085000 ;
      RECT 2.715000  0.085000 2.885000 0.555000 ;
      RECT 3.095000  1.625000 3.345000 2.295000 ;
      RECT 3.095000  2.295000 5.025000 2.465000 ;
      RECT 3.555000  0.085000 3.725000 0.555000 ;
      RECT 3.935000  2.135000 4.185000 2.295000 ;
      RECT 4.395000  0.085000 4.565000 0.555000 ;
      RECT 4.775000  2.135000 5.025000 2.295000 ;
      RECT 5.195000  2.125000 5.445000 2.465000 ;
      RECT 5.235000  0.085000 5.405000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.125000 2.615000 2.295000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.125000 5.375000 2.295000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 2.385000 2.065000 2.680000 2.140000 ;
      RECT 2.385000 2.140000 5.440000 2.280000 ;
      RECT 2.385000 2.280000 2.680000 2.335000 ;
      RECT 5.145000 2.065000 5.440000 2.140000 ;
      RECT 5.145000 2.280000 5.440000 2.335000 ;
  END
END sky130_fd_sc_hd__nor3_4
MACRO sky130_fd_sc_hd__nor3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475000 0.995000 1.815000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.995000 1.305000 1.615000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.995000 2.335000 1.615000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  0.716500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.605000 0.655000 ;
        RECT 0.085000 0.655000 1.445000 0.825000 ;
        RECT 0.085000 0.825000 0.255000 1.445000 ;
        RECT 0.085000 1.445000 0.545000 2.455000 ;
        RECT 1.275000 0.310000 1.445000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.425000  1.075000 0.885000 1.245000 ;
      RECT 0.715000  1.245000 0.885000 1.785000 ;
      RECT 0.715000  1.785000 2.675000 1.955000 ;
      RECT 0.775000  0.085000 1.105000 0.485000 ;
      RECT 1.615000  0.085000 1.945000 0.825000 ;
      RECT 1.615000  2.125000 1.945000 2.635000 ;
      RECT 2.180000  0.405000 2.350000 0.655000 ;
      RECT 2.180000  0.655000 2.675000 0.825000 ;
      RECT 2.505000  0.825000 2.675000 1.785000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__nor3b_1
MACRO sky130_fd_sc_hd__nor3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.965000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135000 1.075000 2.640000 1.285000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.030000 1.075000 4.515000 1.285000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  0.796500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 3.105000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.775000 0.255000 3.105000 0.725000 ;
        RECT 2.815000 0.905000 3.065000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 2.085000 1.625000 ;
      RECT 0.090000  1.625000 0.405000 2.465000 ;
      RECT 0.575000  1.795000 0.825000 2.635000 ;
      RECT 0.995000  1.625000 1.245000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.415000  1.795000 1.665000 2.295000 ;
      RECT 1.415000  2.295000 3.480000 2.465000 ;
      RECT 1.835000  1.625000 2.085000 2.125000 ;
      RECT 1.875000  0.085000 2.605000 0.555000 ;
      RECT 2.375000  1.455000 2.645000 2.295000 ;
      RECT 3.235000  1.075000 3.860000 1.285000 ;
      RECT 3.235000  1.455000 3.480000 2.295000 ;
      RECT 3.275000  0.085000 3.480000 0.895000 ;
      RECT 3.690000  0.380000 4.045000 0.905000 ;
      RECT 3.690000  0.905000 3.860000 1.075000 ;
      RECT 3.690000  1.285000 3.860000 1.455000 ;
      RECT 3.690000  1.455000 4.045000 1.870000 ;
      RECT 4.215000  0.085000 4.505000 0.825000 ;
      RECT 4.215000  1.540000 4.465000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__nor3b_2
MACRO sky130_fd_sc_hd__nor3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 1.075000 2.690000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035000 1.075000 4.300000 1.285000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.445000 1.285000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  1.593000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 0.255000 1.285000 0.725000 ;
        RECT 0.955000 0.725000 6.760000 0.905000 ;
        RECT 1.795000 0.255000 2.125000 0.725000 ;
        RECT 3.155000 0.255000 3.485000 0.725000 ;
        RECT 3.995000 0.255000 4.325000 0.725000 ;
        RECT 4.835000 0.255000 5.165000 0.725000 ;
        RECT 4.875000 1.455000 6.760000 1.625000 ;
        RECT 4.875000 1.625000 5.125000 2.125000 ;
        RECT 5.675000 0.255000 6.005000 0.725000 ;
        RECT 5.715000 1.625000 5.965000 2.125000 ;
        RECT 6.420000 0.905000 6.760000 1.455000 ;
        RECT 6.515000 0.315000 6.760000 0.725000 ;
        RECT 6.555000 1.625000 6.760000 2.415000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.090000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.110000  0.255000 0.445000 0.735000 ;
      RECT 0.110000  0.735000 0.785000 0.905000 ;
      RECT 0.110000  1.455000 4.705000 1.625000 ;
      RECT 0.110000  1.625000 0.405000 2.465000 ;
      RECT 0.575000  1.795000 0.825000 2.635000 ;
      RECT 0.615000  0.085000 0.785000 0.555000 ;
      RECT 0.615000  0.905000 0.785000 1.455000 ;
      RECT 0.995000  1.795000 4.285000 1.965000 ;
      RECT 0.995000  1.965000 1.245000 2.465000 ;
      RECT 1.415000  2.135000 1.665000 2.635000 ;
      RECT 1.455000  0.085000 1.625000 0.555000 ;
      RECT 1.835000  1.965000 2.085000 2.465000 ;
      RECT 2.255000  2.135000 2.505000 2.635000 ;
      RECT 2.295000  0.085000 2.985000 0.555000 ;
      RECT 2.775000  2.135000 3.025000 2.295000 ;
      RECT 2.775000  2.295000 6.385000 2.465000 ;
      RECT 3.195000  1.965000 3.445000 2.125000 ;
      RECT 3.615000  2.135000 3.865000 2.295000 ;
      RECT 3.655000  0.085000 3.825000 0.555000 ;
      RECT 4.035000  1.965000 4.285000 2.125000 ;
      RECT 4.455000  1.795000 4.705000 2.295000 ;
      RECT 4.495000  0.085000 4.665000 0.555000 ;
      RECT 4.535000  1.075000 6.125000 1.285000 ;
      RECT 4.535000  1.285000 4.705000 1.455000 ;
      RECT 5.295000  1.795000 5.545000 2.295000 ;
      RECT 5.335000  0.085000 5.505000 0.555000 ;
      RECT 6.135000  1.795000 6.385000 2.295000 ;
      RECT 6.175000  0.085000 6.345000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
END sky130_fd_sc_hd__nor3b_4
MACRO sky130_fd_sc_hd__nor4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 0.655000 2.215000 1.665000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.245000 1.075000 1.695000 1.245000 ;
        RECT 1.455000 1.245000 1.695000 2.450000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.845000 0.995000 1.075000 1.415000 ;
        RECT 0.845000 1.415000 1.285000 1.615000 ;
        RECT 1.030000 1.615000 1.285000 2.450000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.745000 0.335000 1.325000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.672750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.495000 0.675000 1.665000 ;
        RECT 0.090000 1.665000 0.425000 2.450000 ;
        RECT 0.505000 0.645000 0.860000 0.655000 ;
        RECT 0.505000 0.655000 1.705000 0.825000 ;
        RECT 0.505000 0.825000 0.675000 1.495000 ;
        RECT 0.595000 0.385000 0.860000 0.645000 ;
        RECT 1.535000 0.385000 1.705000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.575000 ;
      RECT 1.035000  0.085000 1.365000 0.485000 ;
      RECT 1.875000  0.085000 2.205000 0.485000 ;
      RECT 1.955000  1.835000 2.215000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4_1
MACRO sky130_fd_sc_hd__nor4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.200000 1.075000 0.965000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135000 1.075000 1.940000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.210000 1.075000 3.105000 1.285000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.340000 1.075000 3.925000 1.285000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.972000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 4.515000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.775000 0.255000 3.105000 0.725000 ;
        RECT 3.615000 0.255000 3.945000 0.725000 ;
        RECT 3.655000 1.455000 4.515000 1.625000 ;
        RECT 3.655000 1.625000 3.905000 2.125000 ;
        RECT 4.180000 0.905000 4.515000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.150000  1.455000 2.085000 1.625000 ;
      RECT 0.150000  1.625000 0.405000 2.465000 ;
      RECT 0.575000  1.795000 0.825000 2.635000 ;
      RECT 0.995000  1.625000 1.245000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.415000  1.795000 1.665000 2.295000 ;
      RECT 1.415000  2.295000 3.065000 2.465000 ;
      RECT 1.835000  1.625000 2.085000 2.125000 ;
      RECT 1.875000  0.085000 2.605000 0.555000 ;
      RECT 2.395000  1.455000 3.485000 1.625000 ;
      RECT 2.395000  1.625000 2.645000 2.125000 ;
      RECT 2.815000  1.795000 3.065000 2.295000 ;
      RECT 3.235000  1.625000 3.485000 2.295000 ;
      RECT 3.235000  2.295000 4.325000 2.465000 ;
      RECT 3.275000  0.085000 3.445000 0.555000 ;
      RECT 4.075000  1.795000 4.325000 2.295000 ;
      RECT 4.115000  0.085000 4.405000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4_2
MACRO sky130_fd_sc_hd__nor4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.180000 1.075000 1.825000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095000 1.075000 4.070000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.295000 1.075000 5.705000 1.285000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.875000 1.075000 7.295000 1.285000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.944000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 7.735000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.215000 0.255000 2.545000 0.725000 ;
        RECT 3.055000 0.255000 3.385000 0.725000 ;
        RECT 4.415000 0.255000 4.745000 0.725000 ;
        RECT 5.255000 0.255000 5.585000 0.725000 ;
        RECT 6.095000 0.255000 6.425000 0.725000 ;
        RECT 6.135000 1.455000 7.735000 1.625000 ;
        RECT 6.135000 1.625000 6.385000 2.125000 ;
        RECT 6.935000 0.255000 7.265000 0.725000 ;
        RECT 6.975000 1.625000 7.225000 2.125000 ;
        RECT 7.465000 0.905000 7.735000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 2.085000 1.625000 ;
      RECT 0.090000  1.625000 0.405000 2.465000 ;
      RECT 0.575000  1.795000 0.825000 2.635000 ;
      RECT 0.995000  1.625000 1.245000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.415000  1.795000 1.665000 2.635000 ;
      RECT 1.835000  1.625000 2.085000 2.295000 ;
      RECT 1.835000  2.295000 3.820000 2.465000 ;
      RECT 1.875000  0.085000 2.045000 0.555000 ;
      RECT 2.255000  1.455000 5.545000 1.625000 ;
      RECT 2.255000  1.625000 2.505000 2.125000 ;
      RECT 2.675000  1.795000 2.925000 2.295000 ;
      RECT 2.715000  0.085000 2.885000 0.555000 ;
      RECT 3.095000  1.625000 3.345000 2.125000 ;
      RECT 3.515000  1.795000 3.820000 2.295000 ;
      RECT 3.555000  0.085000 4.245000 0.555000 ;
      RECT 4.005000  1.795000 4.285000 2.295000 ;
      RECT 4.005000  2.295000 7.645000 2.465000 ;
      RECT 4.455000  1.625000 4.705000 2.125000 ;
      RECT 4.875000  1.795000 5.125000 2.295000 ;
      RECT 4.915000  0.085000 5.085000 0.555000 ;
      RECT 5.295000  1.625000 5.545000 2.125000 ;
      RECT 5.715000  1.795000 5.965000 2.295000 ;
      RECT 5.755000  0.085000 5.925000 0.555000 ;
      RECT 6.555000  1.795000 6.805000 2.295000 ;
      RECT 6.595000  0.085000 6.765000 0.555000 ;
      RECT 7.395000  1.795000 7.645000 2.295000 ;
      RECT 7.435000  0.085000 7.605000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4_4
MACRO sky130_fd_sc_hd__nor4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 0.995000 2.275000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.995000 1.785000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 0.995000 1.285000 1.615000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 0.995000 2.795000 1.615000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.871000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.655000 1.925000 0.825000 ;
        RECT 0.085000 0.825000 0.345000 2.450000 ;
        RECT 0.855000 0.300000 1.055000 0.655000 ;
        RECT 1.725000 0.310000 1.925000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.355000  0.085000 0.685000 0.480000 ;
      RECT 0.525000  0.995000 0.745000 1.795000 ;
      RECT 0.525000  1.795000 3.135000 2.005000 ;
      RECT 1.225000  0.085000 1.555000 0.485000 ;
      RECT 2.095000  0.085000 2.425000 0.825000 ;
      RECT 2.095000  2.185000 2.425000 2.635000 ;
      RECT 2.660000  0.405000 2.830000 0.655000 ;
      RECT 2.660000  0.655000 3.135000 0.825000 ;
      RECT 2.965000  0.825000 3.135000 1.795000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4b_1
MACRO sky130_fd_sc_hd__nor4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.075000 1.240000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.420000 1.075000 2.635000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.815000 1.075000 3.535000 1.285000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.805000 1.075000 5.435000 1.285000 ;
        RECT 5.185000 1.285000 5.435000 1.955000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.972000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.845000 0.725000 ;
        RECT 0.515000 0.725000 3.920000 0.905000 ;
        RECT 1.355000 0.255000 1.685000 0.725000 ;
        RECT 2.750000 0.255000 3.080000 0.725000 ;
        RECT 3.590000 0.255000 3.920000 0.725000 ;
        RECT 3.630000 1.455000 4.035000 1.625000 ;
        RECT 3.630000 1.625000 3.880000 2.125000 ;
        RECT 3.715000 0.905000 3.920000 1.075000 ;
        RECT 3.715000 1.075000 4.035000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.905000 ;
      RECT 0.085000  1.455000 2.105000 1.625000 ;
      RECT 0.085000  1.625000 0.425000 2.465000 ;
      RECT 0.595000  1.795000 0.805000 2.635000 ;
      RECT 0.975000  1.625000 1.225000 2.465000 ;
      RECT 1.015000  0.085000 1.185000 0.555000 ;
      RECT 1.395000  1.795000 1.605000 2.295000 ;
      RECT 1.395000  2.295000 3.040000 2.465000 ;
      RECT 1.775000  1.625000 2.105000 2.125000 ;
      RECT 1.855000  0.085000 2.580000 0.555000 ;
      RECT 2.275000  1.455000 3.460000 1.625000 ;
      RECT 2.275000  1.625000 2.660000 2.125000 ;
      RECT 2.830000  1.795000 3.040000 2.295000 ;
      RECT 3.210000  1.625000 3.460000 2.295000 ;
      RECT 3.210000  2.295000 4.295000 2.465000 ;
      RECT 3.250000  0.085000 3.420000 0.555000 ;
      RECT 4.050000  1.795000 4.295000 2.295000 ;
      RECT 4.090000  0.085000 4.295000 0.895000 ;
      RECT 4.320000  1.075000 4.635000 1.245000 ;
      RECT 4.465000  0.380000 4.820000 0.905000 ;
      RECT 4.465000  0.905000 4.635000 1.075000 ;
      RECT 4.465000  1.245000 4.635000 2.035000 ;
      RECT 4.465000  2.035000 4.820000 2.450000 ;
      RECT 4.990000  0.085000 5.240000 0.825000 ;
      RECT 4.990000  2.135000 5.240000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4b_2
MACRO sky130_fd_sc_hd__nor4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.395000 1.075000 1.805000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.075000 3.750000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.985000 1.075000 5.685000 1.285000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.810000 1.075000 8.655000 1.285000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.944000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.845000 0.725000 ;
        RECT 0.515000 0.725000 7.245000 0.905000 ;
        RECT 1.355000 0.255000 1.685000 0.725000 ;
        RECT 2.195000 0.255000 2.525000 0.725000 ;
        RECT 3.035000 0.255000 3.365000 0.725000 ;
        RECT 4.395000 0.255000 4.725000 0.725000 ;
        RECT 5.235000 0.255000 5.565000 0.725000 ;
        RECT 6.075000 0.255000 6.405000 0.725000 ;
        RECT 6.115000 0.905000 6.465000 1.455000 ;
        RECT 6.115000 1.455000 7.205000 1.625000 ;
        RECT 6.115000 1.625000 6.365000 2.125000 ;
        RECT 6.915000 0.255000 7.245000 0.725000 ;
        RECT 6.955000 1.625000 7.205000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.930000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.095000  1.455000 2.065000 1.625000 ;
      RECT 0.095000  1.625000 0.425000 2.465000 ;
      RECT 0.175000  0.085000 0.345000 0.895000 ;
      RECT 0.595000  1.795000 0.805000 2.635000 ;
      RECT 0.975000  1.625000 1.225000 2.465000 ;
      RECT 1.015000  0.085000 1.185000 0.555000 ;
      RECT 1.395000  1.795000 1.645000 2.635000 ;
      RECT 1.815000  1.625000 2.065000 2.295000 ;
      RECT 1.815000  2.295000 3.745000 2.465000 ;
      RECT 1.855000  0.085000 2.025000 0.555000 ;
      RECT 2.235000  1.455000 5.525000 1.625000 ;
      RECT 2.235000  1.625000 2.485000 2.125000 ;
      RECT 2.655000  1.795000 2.905000 2.295000 ;
      RECT 2.695000  0.085000 2.865000 0.555000 ;
      RECT 3.075000  1.625000 3.325000 2.125000 ;
      RECT 3.495000  1.795000 3.745000 2.295000 ;
      RECT 3.535000  0.085000 4.225000 0.555000 ;
      RECT 4.015000  1.795000 4.265000 2.295000 ;
      RECT 4.015000  2.295000 7.625000 2.465000 ;
      RECT 4.435000  1.625000 4.685000 2.125000 ;
      RECT 4.855000  1.795000 5.105000 2.295000 ;
      RECT 4.895000  0.085000 5.065000 0.555000 ;
      RECT 5.275000  1.625000 5.525000 2.125000 ;
      RECT 5.695000  1.455000 5.945000 2.295000 ;
      RECT 5.735000  0.085000 5.905000 0.555000 ;
      RECT 6.535000  1.795000 6.785000 2.295000 ;
      RECT 6.575000  0.085000 6.745000 0.555000 ;
      RECT 6.635000  1.075000 7.640000 1.285000 ;
      RECT 7.375000  1.795000 7.625000 2.295000 ;
      RECT 7.415000  0.085000 7.585000 0.555000 ;
      RECT 7.470000  0.735000 8.185000 0.905000 ;
      RECT 7.470000  0.905000 7.640000 1.075000 ;
      RECT 7.470000  1.285000 7.640000 1.455000 ;
      RECT 7.470000  1.455000 8.185000 1.625000 ;
      RECT 7.810000  0.255000 8.185000 0.735000 ;
      RECT 7.850000  1.625000 8.185000 2.465000 ;
      RECT 8.355000  0.085000 8.585000 0.905000 ;
      RECT 8.355000  1.455000 8.585000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4b_4
MACRO sky130_fd_sc_hd__nor4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.115000 0.995000 3.595000 1.275000 ;
        RECT 3.295000 1.275000 3.595000 1.705000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615000 0.995000 2.945000 1.445000 ;
        RECT 2.615000 1.445000 3.085000 1.630000 ;
        RECT 2.825000 1.630000 3.085000 2.410000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.995000 0.780000 1.695000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.995000 1.240000 1.325000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.606900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.470000 1.955000 2.055000 2.125000 ;
        RECT 1.855000 0.655000 3.085000 0.825000 ;
        RECT 1.855000 0.825000 2.055000 1.955000 ;
        RECT 2.015000 0.300000 2.215000 0.655000 ;
        RECT 2.885000 0.310000 3.085000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.450000 0.405000 0.825000 ;
      RECT 0.085000  0.825000 0.260000 1.885000 ;
      RECT 0.085000  1.885000 1.205000 2.070000 ;
      RECT 0.085000  2.070000 0.345000 2.455000 ;
      RECT 0.515000  2.240000 0.845000 2.635000 ;
      RECT 0.655000  0.085000 0.825000 0.825000 ;
      RECT 0.995000  1.525000 1.590000 1.715000 ;
      RECT 1.035000  2.070000 1.205000 2.295000 ;
      RECT 1.035000  2.295000 2.395000 2.465000 ;
      RECT 1.075000  0.450000 1.245000 0.655000 ;
      RECT 1.075000  0.655000 1.590000 0.825000 ;
      RECT 1.410000  0.825000 1.590000 0.995000 ;
      RECT 1.410000  0.995000 1.685000 1.325000 ;
      RECT 1.410000  1.325000 1.590000 1.525000 ;
      RECT 1.515000  0.085000 1.845000 0.480000 ;
      RECT 2.225000  0.995000 2.395000 2.295000 ;
      RECT 2.385000  0.085000 2.715000 0.485000 ;
      RECT 3.255000  0.085000 3.585000 0.825000 ;
      RECT 3.255000  1.875000 3.585000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4bb_1
MACRO sky130_fd_sc_hd__nor4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.130000 1.075000 5.895000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165000 1.075000 4.960000 1.275000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.995000 1.235000 1.325000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.780000 1.695000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.972000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.060000 0.255000 2.390000 0.725000 ;
        RECT 2.060000 0.725000 5.450000 0.905000 ;
        RECT 2.900000 0.255000 3.230000 0.725000 ;
        RECT 2.900000 1.445000 3.995000 1.705000 ;
        RECT 3.575000 0.905000 3.995000 1.445000 ;
        RECT 4.280000 0.255000 4.610000 0.725000 ;
        RECT 5.120000 0.255000 5.450000 0.725000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.450000 0.465000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.885000 ;
      RECT 0.085000  1.885000 1.915000 2.055000 ;
      RECT 0.085000  2.055000 0.345000 2.455000 ;
      RECT 0.515000  2.240000 0.845000 2.635000 ;
      RECT 0.635000  0.085000 0.805000 0.825000 ;
      RECT 0.995000  1.525000 1.575000 1.715000 ;
      RECT 1.055000  0.450000 1.250000 0.655000 ;
      RECT 1.055000  0.655000 1.575000 0.825000 ;
      RECT 1.405000  0.825000 1.575000 1.075000 ;
      RECT 1.405000  1.075000 2.390000 1.245000 ;
      RECT 1.405000  1.245000 1.575000 1.525000 ;
      RECT 1.560000  0.085000 1.890000 0.480000 ;
      RECT 1.640000  2.225000 1.970000 2.295000 ;
      RECT 1.640000  2.295000 3.650000 2.465000 ;
      RECT 1.745000  1.415000 2.730000 1.585000 ;
      RECT 1.745000  1.585000 1.915000 1.885000 ;
      RECT 2.140000  1.795000 2.310000 1.875000 ;
      RECT 2.140000  1.875000 4.610000 2.045000 ;
      RECT 2.140000  2.045000 2.310000 2.125000 ;
      RECT 2.480000  2.215000 3.650000 2.295000 ;
      RECT 2.560000  0.085000 2.730000 0.555000 ;
      RECT 2.560000  1.075000 3.405000 1.275000 ;
      RECT 2.560000  1.275000 2.730000 1.415000 ;
      RECT 3.400000  0.085000 4.110000 0.555000 ;
      RECT 3.860000  2.215000 4.990000 2.465000 ;
      RECT 4.320000  1.455000 4.610000 1.875000 ;
      RECT 4.780000  0.085000 4.950000 0.555000 ;
      RECT 4.780000  1.455000 5.870000 1.625000 ;
      RECT 4.780000  1.625000 4.990000 2.215000 ;
      RECT 5.160000  1.795000 5.370000 2.635000 ;
      RECT 5.540000  1.625000 5.870000 2.465000 ;
      RECT 5.620000  0.085000 5.895000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4bb_2
MACRO sky130_fd_sc_hd__nor4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.375000 1.075000 9.110000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.150000 1.075000 7.105000 1.285000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.445000 1.365000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 1.075000 1.295000 1.325000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.944000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.840000 1.415000 3.185000 1.705000 ;
        RECT 1.935000 0.255000 2.265000 0.725000 ;
        RECT 1.935000 0.725000 8.665000 0.905000 ;
        RECT 2.775000 0.255000 3.105000 0.725000 ;
        RECT 3.015000 0.905000 3.185000 1.415000 ;
        RECT 3.615000 0.255000 3.945000 0.725000 ;
        RECT 4.455000 0.255000 4.785000 0.725000 ;
        RECT 5.815000 0.255000 6.145000 0.725000 ;
        RECT 6.655000 0.255000 6.985000 0.725000 ;
        RECT 7.495000 0.255000 7.825000 0.725000 ;
        RECT 8.335000 0.255000 8.665000 0.725000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.085000  0.255000 0.445000 0.725000 ;
      RECT 0.085000  0.725000 0.785000 0.895000 ;
      RECT 0.085000  1.535000 0.785000 1.875000 ;
      RECT 0.085000  1.875000 3.525000 2.045000 ;
      RECT 0.085000  2.045000 0.365000 2.465000 ;
      RECT 0.535000  2.215000 0.865000 2.635000 ;
      RECT 0.615000  0.085000 0.785000 0.555000 ;
      RECT 0.615000  0.895000 0.785000 1.535000 ;
      RECT 0.955000  0.255000 1.285000 0.735000 ;
      RECT 0.955000  0.735000 1.635000 0.905000 ;
      RECT 0.955000  1.535000 1.635000 1.705000 ;
      RECT 1.465000  0.905000 1.635000 1.075000 ;
      RECT 1.465000  1.075000 2.845000 1.245000 ;
      RECT 1.465000  1.245000 1.635000 1.535000 ;
      RECT 1.515000  2.215000 3.525000 2.295000 ;
      RECT 1.515000  2.295000 5.195000 2.465000 ;
      RECT 1.595000  0.085000 1.765000 0.555000 ;
      RECT 2.435000  0.085000 2.605000 0.555000 ;
      RECT 3.275000  0.085000 3.445000 0.555000 ;
      RECT 3.355000  1.075000 4.905000 1.285000 ;
      RECT 3.355000  1.285000 3.525000 1.875000 ;
      RECT 3.695000  1.455000 6.945000 1.625000 ;
      RECT 3.695000  1.625000 3.905000 2.125000 ;
      RECT 4.075000  1.795000 4.325000 2.295000 ;
      RECT 4.115000  0.085000 4.285000 0.555000 ;
      RECT 4.495000  1.625000 4.745000 2.125000 ;
      RECT 4.915000  1.795000 5.195000 2.295000 ;
      RECT 4.955000  0.085000 5.645000 0.555000 ;
      RECT 5.380000  1.795000 5.685000 2.295000 ;
      RECT 5.380000  2.295000 7.365000 2.465000 ;
      RECT 5.855000  1.625000 6.105000 2.125000 ;
      RECT 6.275000  1.795000 6.525000 2.295000 ;
      RECT 6.315000  0.085000 6.485000 0.555000 ;
      RECT 6.695000  1.625000 6.945000 2.125000 ;
      RECT 7.115000  1.455000 9.110000 1.625000 ;
      RECT 7.115000  1.625000 7.365000 2.295000 ;
      RECT 7.155000  0.085000 7.325000 0.555000 ;
      RECT 7.535000  1.795000 7.785000 2.635000 ;
      RECT 7.955000  1.625000 8.205000 2.465000 ;
      RECT 7.995000  0.085000 8.165000 0.555000 ;
      RECT 8.375000  1.795000 8.625000 2.635000 ;
      RECT 8.795000  1.625000 9.110000 2.465000 ;
      RECT 8.835000  0.085000 9.110000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4bb_4
MACRO sky130_fd_sc_hd__o2bb2a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.770000 1.075000 1.220000 1.275000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 0.380000 1.290000 0.735000 ;
        RECT 1.070000 0.735000 1.565000 0.905000 ;
        RECT 1.390000 0.905000 1.565000 1.100000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.250000 1.075000 3.595000 1.645000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.520000 1.075000 3.080000 1.325000 ;
        RECT 2.905000 1.325000 3.080000 2.425000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.425000 0.825000 ;
        RECT 0.085000 0.825000 0.260000 1.795000 ;
        RECT 0.085000 1.795000 0.345000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.430000  0.995000 0.600000 1.445000 ;
      RECT 0.430000  1.445000 0.825000 1.615000 ;
      RECT 0.515000  2.235000 0.845000 2.635000 ;
      RECT 0.620000  0.085000 0.790000 0.750000 ;
      RECT 0.655000  1.615000 0.825000 1.885000 ;
      RECT 0.655000  1.885000 2.735000 2.055000 ;
      RECT 0.995000  1.495000 2.010000 1.715000 ;
      RECT 1.460000  0.395000 1.905000 0.565000 ;
      RECT 1.715000  2.235000 2.115000 2.635000 ;
      RECT 1.735000  0.565000 1.905000 1.355000 ;
      RECT 1.735000  1.355000 2.010000 1.495000 ;
      RECT 2.075000  0.320000 2.325000 0.690000 ;
      RECT 2.155000  0.690000 2.325000 1.075000 ;
      RECT 2.155000  1.075000 2.350000 1.245000 ;
      RECT 2.180000  1.245000 2.350000 1.495000 ;
      RECT 2.180000  1.495000 2.735000 1.885000 ;
      RECT 2.405000  2.055000 2.735000 2.290000 ;
      RECT 2.495000  0.320000 2.745000 0.725000 ;
      RECT 2.495000  0.725000 3.595000 0.905000 ;
      RECT 2.915000  0.085000 3.085000 0.555000 ;
      RECT 3.250000  1.815000 3.595000 2.635000 ;
      RECT 3.255000  0.320000 3.595000 0.725000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o2bb2a_1
MACRO sky130_fd_sc_hd__o2bb2a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.215000 1.075000 1.685000 1.275000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 0.380000 1.735000 0.735000 ;
        RECT 1.515000 0.735000 2.020000 0.770000 ;
        RECT 1.515000 0.770000 2.025000 0.905000 ;
        RECT 1.855000 0.905000 2.025000 1.100000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.700000 1.075000 4.045000 1.645000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.075000 3.525000 1.325000 ;
        RECT 3.355000 1.325000 3.525000 2.425000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.870000 0.825000 ;
        RECT 0.535000 0.825000 0.705000 1.795000 ;
        RECT 0.535000 1.795000 0.790000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.135000 -0.085000 0.305000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.110000  0.085000 0.365000 0.910000 ;
      RECT 0.110000  1.410000 0.365000 2.635000 ;
      RECT 0.875000  0.995000 1.045000 1.445000 ;
      RECT 0.875000  1.445000 1.270000 1.615000 ;
      RECT 0.960000  2.235000 1.290000 2.635000 ;
      RECT 1.065000  0.085000 1.235000 0.750000 ;
      RECT 1.100000  1.615000 1.270000 1.885000 ;
      RECT 1.100000  1.885000 3.185000 2.055000 ;
      RECT 1.440000  1.495000 2.460000 1.715000 ;
      RECT 1.905000  0.395000 2.365000 0.565000 ;
      RECT 2.160000  2.235000 2.565000 2.635000 ;
      RECT 2.195000  0.565000 2.365000 1.355000 ;
      RECT 2.195000  1.355000 2.460000 1.495000 ;
      RECT 2.535000  0.320000 2.780000 0.690000 ;
      RECT 2.610000  0.690000 2.780000 1.075000 ;
      RECT 2.610000  1.075000 2.800000 1.245000 ;
      RECT 2.630000  1.245000 2.800000 1.495000 ;
      RECT 2.630000  1.495000 3.185000 1.885000 ;
      RECT 2.835000  2.055000 3.185000 2.425000 ;
      RECT 2.955000  0.320000 3.185000 0.725000 ;
      RECT 2.955000  0.725000 4.045000 0.905000 ;
      RECT 3.375000  0.085000 3.545000 0.555000 ;
      RECT 3.715000  0.320000 4.045000 0.725000 ;
      RECT 3.730000  1.815000 4.045000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__o2bb2a_2
MACRO sky130_fd_sc_hd__o2bb2a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 1.075000 3.645000 1.445000 ;
        RECT 3.315000 1.445000 4.965000 1.615000 ;
        RECT 4.605000 1.075000 4.965000 1.445000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 1.075000 4.435000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.575000 1.445000 ;
        RECT 0.085000 1.445000 1.895000 1.615000 ;
        RECT 1.565000 1.075000 1.895000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 1.075000 1.345000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235000 0.275000 5.565000 0.725000 ;
        RECT 5.235000 0.725000 6.910000 0.905000 ;
        RECT 5.275000 1.785000 6.365000 1.955000 ;
        RECT 5.275000 1.955000 5.525000 2.465000 ;
        RECT 6.075000 0.275000 6.405000 0.725000 ;
        RECT 6.115000 1.415000 6.910000 1.655000 ;
        RECT 6.115000 1.655000 6.365000 1.785000 ;
        RECT 6.115000 1.955000 6.365000 2.465000 ;
        RECT 6.605000 0.905000 6.910000 1.415000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.095000  0.255000 0.425000 0.725000 ;
      RECT 0.095000  0.725000 1.265000 0.735000 ;
      RECT 0.095000  0.735000 2.025000 0.905000 ;
      RECT 0.140000  1.795000 0.345000 2.635000 ;
      RECT 0.555000  1.785000 0.805000 2.295000 ;
      RECT 0.555000  2.295000 1.645000 2.465000 ;
      RECT 0.595000  0.085000 0.765000 0.555000 ;
      RECT 0.935000  0.255000 1.265000 0.725000 ;
      RECT 0.975000  1.785000 2.615000 1.955000 ;
      RECT 0.975000  1.955000 1.225000 2.125000 ;
      RECT 1.395000  2.125000 1.645000 2.295000 ;
      RECT 1.435000  0.085000 1.605000 0.555000 ;
      RECT 1.775000  0.255000 2.945000 0.475000 ;
      RECT 1.775000  0.475000 2.025000 0.735000 ;
      RECT 1.815000  2.125000 2.065000 2.635000 ;
      RECT 2.065000  1.075000 2.445000 1.415000 ;
      RECT 2.065000  1.415000 2.615000 1.785000 ;
      RECT 2.195000  0.645000 2.525000 0.815000 ;
      RECT 2.195000  0.815000 2.445000 1.075000 ;
      RECT 2.235000  1.955000 2.615000 1.965000 ;
      RECT 2.235000  1.965000 2.525000 2.465000 ;
      RECT 2.615000  1.075000 3.145000 1.245000 ;
      RECT 2.695000  2.135000 3.425000 2.635000 ;
      RECT 2.955000  0.725000 4.305000 0.905000 ;
      RECT 2.955000  0.905000 3.145000 1.075000 ;
      RECT 2.955000  1.245000 3.145000 1.785000 ;
      RECT 2.955000  1.785000 4.685000 1.965000 ;
      RECT 3.215000  0.085000 3.385000 0.555000 ;
      RECT 3.555000  0.305000 4.725000 0.475000 ;
      RECT 3.595000  1.965000 3.845000 2.125000 ;
      RECT 3.975000  0.645000 4.305000 0.725000 ;
      RECT 4.015000  2.135000 4.265000 2.635000 ;
      RECT 4.435000  1.965000 4.685000 2.465000 ;
      RECT 4.475000  0.475000 4.725000 0.895000 ;
      RECT 4.855000  1.795000 5.105000 2.635000 ;
      RECT 4.895000  0.085000 5.065000 0.895000 ;
      RECT 5.165000  1.075000 6.435000 1.245000 ;
      RECT 5.165000  1.245000 5.455000 1.615000 ;
      RECT 5.695000  2.165000 5.945000 2.635000 ;
      RECT 5.735000  0.085000 5.905000 0.555000 ;
      RECT 6.535000  1.825000 6.785000 2.635000 ;
      RECT 6.575000  0.085000 6.745000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  1.445000 2.615000 1.615000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.225000  1.445000 5.395000 1.615000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
    LAYER met1 ;
      RECT 2.385000 1.415000 2.675000 1.460000 ;
      RECT 2.385000 1.460000 5.455000 1.600000 ;
      RECT 2.385000 1.600000 2.675000 1.645000 ;
      RECT 5.165000 1.415000 5.455000 1.460000 ;
      RECT 5.165000 1.600000 5.455000 1.645000 ;
  END
END sky130_fd_sc_hd__o2bb2a_4
MACRO sky130_fd_sc_hd__o2bb2ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.435000 1.285000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.280000 0.825000 0.995000 ;
        RECT 0.605000 0.995000 1.000000 1.325000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 1.075000 3.135000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.030000 1.075000 2.615000 1.325000 ;
        RECT 2.445000 1.325000 2.615000 2.425000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.560000 0.430000 1.810000 0.790000 ;
        RECT 1.640000 0.790000 1.810000 1.495000 ;
        RECT 1.640000 1.495000 2.270000 1.665000 ;
        RECT 1.940000 1.665000 2.270000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.815000 ;
      RECT 0.150000  1.455000 0.400000 2.635000 ;
      RECT 0.570000  1.495000 1.340000 1.665000 ;
      RECT 0.570000  1.665000 0.820000 2.465000 ;
      RECT 0.990000  1.835000 1.770000 2.635000 ;
      RECT 1.000000  0.280000 1.340000 0.825000 ;
      RECT 1.170000  0.825000 1.340000 0.995000 ;
      RECT 1.170000  0.995000 1.470000 1.325000 ;
      RECT 1.170000  1.325000 1.340000 1.495000 ;
      RECT 1.980000  0.425000 2.270000 0.725000 ;
      RECT 1.980000  0.725000 3.110000 0.905000 ;
      RECT 2.440000  0.085000 2.610000 0.555000 ;
      RECT 2.780000  0.275000 3.110000 0.725000 ;
      RECT 2.820000  1.455000 3.070000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o2bb2ai_1
MACRO sky130_fd_sc_hd__o2bb2ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.625000 1.445000 ;
        RECT 0.090000 1.445000 1.945000 1.615000 ;
        RECT 1.615000 1.075000 1.945000 1.445000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.795000 1.075000 1.400000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.410000 1.075000 3.740000 1.445000 ;
        RECT 3.410000 1.445000 5.435000 1.615000 ;
        RECT 4.730000 1.075000 5.435000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.960000 1.075000 4.500000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.745000 0.645000 3.075000 1.075000 ;
        RECT 2.745000 1.075000 3.215000 1.785000 ;
        RECT 2.745000 1.785000 4.330000 1.955000 ;
        RECT 2.745000 1.955000 3.035000 2.465000 ;
        RECT 4.080000 1.955000 4.330000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.150000  1.795000 0.400000 2.635000 ;
      RECT 0.195000  0.085000 0.365000 0.895000 ;
      RECT 0.535000  0.305000 1.705000 0.475000 ;
      RECT 0.535000  0.475000 0.785000 0.895000 ;
      RECT 0.575000  1.785000 2.285000 1.965000 ;
      RECT 0.575000  1.965000 0.825000 2.465000 ;
      RECT 0.955000  0.645000 1.285000 0.725000 ;
      RECT 0.955000  0.725000 2.285000 0.905000 ;
      RECT 0.995000  2.135000 1.245000 2.635000 ;
      RECT 1.415000  1.965000 1.665000 2.125000 ;
      RECT 1.835000  2.135000 2.575000 2.635000 ;
      RECT 1.875000  0.085000 2.045000 0.555000 ;
      RECT 2.115000  0.905000 2.285000 0.995000 ;
      RECT 2.115000  0.995000 2.575000 1.325000 ;
      RECT 2.115000  1.325000 2.285000 1.785000 ;
      RECT 2.325000  0.255000 3.530000 0.475000 ;
      RECT 2.325000  0.475000 2.575000 0.555000 ;
      RECT 3.205000  2.125000 3.490000 2.635000 ;
      RECT 3.245000  0.475000 3.530000 0.735000 ;
      RECT 3.245000  0.735000 5.210000 0.905000 ;
      RECT 3.660000  2.125000 3.910000 2.295000 ;
      RECT 3.660000  2.295000 4.750000 2.465000 ;
      RECT 3.700000  0.085000 3.870000 0.555000 ;
      RECT 4.040000  0.255000 4.370000 0.725000 ;
      RECT 4.040000  0.725000 5.210000 0.735000 ;
      RECT 4.500000  1.785000 4.750000 2.295000 ;
      RECT 4.540000  0.085000 4.710000 0.555000 ;
      RECT 4.880000  0.255000 5.210000 0.725000 ;
      RECT 4.965000  1.795000 5.170000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__o2bb2ai_2
MACRO sky130_fd_sc_hd__o2bb2ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095000 1.075000 3.505000 1.285000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 1.825000 1.285000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.045000 1.075000 10.005000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.465000 1.075000 7.875000 1.285000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.415000 0.645000 6.155000 0.905000 ;
        RECT 4.425000 1.455000 7.715000 1.625000 ;
        RECT 4.425000 1.625000 4.675000 2.465000 ;
        RECT 5.265000 1.625000 5.515000 2.465000 ;
        RECT 5.875000 0.905000 6.155000 1.455000 ;
        RECT 6.625000 1.625000 6.875000 2.125000 ;
        RECT 7.465000 1.625000 7.715000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.135000 -0.085000 0.305000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.085000  0.645000  1.705000 0.905000 ;
      RECT 0.085000  0.905000  0.255000 1.455000 ;
      RECT 0.085000  1.455000  3.915000 1.625000 ;
      RECT 0.100000  0.255000  2.125000 0.475000 ;
      RECT 0.155000  1.795000  0.405000 2.635000 ;
      RECT 0.575000  1.625000  0.825000 2.465000 ;
      RECT 0.995000  1.795000  1.245000 2.635000 ;
      RECT 1.415000  1.625000  1.665000 2.465000 ;
      RECT 1.835000  1.795000  2.085000 2.635000 ;
      RECT 1.875000  0.475000  2.125000 0.725000 ;
      RECT 1.875000  0.725000  3.805000 0.905000 ;
      RECT 2.255000  1.625000  2.505000 2.465000 ;
      RECT 2.295000  0.085000  2.465000 0.555000 ;
      RECT 2.635000  0.255000  2.965000 0.725000 ;
      RECT 2.675000  1.795000  2.925000 2.635000 ;
      RECT 3.095000  1.625000  3.345000 2.465000 ;
      RECT 3.135000  0.085000  3.305000 0.555000 ;
      RECT 3.475000  0.255000  3.805000 0.725000 ;
      RECT 3.515000  1.795000  4.255000 2.635000 ;
      RECT 3.745000  1.075000  5.705000 1.285000 ;
      RECT 3.745000  1.285000  3.915000 1.455000 ;
      RECT 4.060000  0.255000  6.495000 0.475000 ;
      RECT 4.060000  0.475000  4.245000 0.835000 ;
      RECT 4.845000  1.795000  5.095000 2.635000 ;
      RECT 5.685000  1.795000  5.935000 2.635000 ;
      RECT 6.175000  1.795000  6.455000 2.295000 ;
      RECT 6.175000  2.295000  8.135000 2.465000 ;
      RECT 6.325000  0.475000  6.495000 0.735000 ;
      RECT 6.325000  0.735000  9.855000 0.905000 ;
      RECT 6.665000  0.085000  6.835000 0.555000 ;
      RECT 7.005000  0.255000  7.335000 0.725000 ;
      RECT 7.005000  0.725000  9.855000 0.735000 ;
      RECT 7.045000  1.795000  7.295000 2.295000 ;
      RECT 7.505000  0.085000  7.675000 0.555000 ;
      RECT 7.845000  0.255000  8.175000 0.725000 ;
      RECT 7.885000  1.455000  9.875000 1.625000 ;
      RECT 7.885000  1.625000  8.135000 2.295000 ;
      RECT 8.305000  1.795000  8.555000 2.635000 ;
      RECT 8.345000  0.085000  8.515000 0.555000 ;
      RECT 8.685000  0.255000  9.015000 0.725000 ;
      RECT 8.725000  1.625000  8.975000 2.465000 ;
      RECT 9.145000  1.795000  9.395000 2.635000 ;
      RECT 9.185000  0.085000  9.355000 0.555000 ;
      RECT 9.525000  0.255000  9.855000 0.725000 ;
      RECT 9.565000  1.625000  9.875000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
END sky130_fd_sc_hd__o2bb2ai_4
MACRO sky130_fd_sc_hd__o21a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.345000 1.075000 2.675000 1.275000 ;
        RECT 2.445000 1.275000 2.675000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.705000 1.075000 2.035000 1.095000 ;
        RECT 1.705000 1.095000 2.155000 1.275000 ;
        RECT 1.940000 1.275000 2.155000 2.390000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.075000 1.535000 1.305000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.425000 1.030000 ;
        RECT 0.085000 1.030000 0.365000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.535000  1.860000 1.245000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.545000 ;
      RECT 0.595000  0.715000 1.305000 0.905000 ;
      RECT 0.595000  0.905000 0.880000 1.475000 ;
      RECT 0.595000  1.475000 1.745000 1.690000 ;
      RECT 1.005000  0.255000 1.365000 0.520000 ;
      RECT 1.005000  0.520000 1.360000 0.525000 ;
      RECT 1.005000  0.525000 1.355000 0.535000 ;
      RECT 1.005000  0.535000 1.350000 0.540000 ;
      RECT 1.005000  0.540000 1.345000 0.550000 ;
      RECT 1.005000  0.550000 1.340000 0.555000 ;
      RECT 1.005000  0.555000 1.330000 0.565000 ;
      RECT 1.005000  0.565000 1.320000 0.575000 ;
      RECT 1.005000  0.575000 1.305000 0.715000 ;
      RECT 1.415000  1.690000 1.745000 2.465000 ;
      RECT 1.495000  0.635000 1.825000 0.715000 ;
      RECT 1.495000  0.715000 2.675000 0.905000 ;
      RECT 1.995000  0.085000 2.165000 0.545000 ;
      RECT 2.335000  0.255000 2.675000 0.715000 ;
      RECT 2.335000  1.915000 2.665000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__o21a_1
MACRO sky130_fd_sc_hd__o21a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865000 0.995000 3.125000 1.450000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025000 1.025000 2.610000 1.400000 ;
        RECT 2.405000 1.400000 2.610000 1.985000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445000 1.010000 1.855000 1.615000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.530000 0.255000 0.775000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  1.635000 0.345000 2.635000 ;
      RECT 0.105000  0.085000 0.345000 0.885000 ;
      RECT 0.945000  0.085000 1.275000 0.465000 ;
      RECT 0.945000  0.635000 1.795000 0.840000 ;
      RECT 0.945000  0.840000 1.275000 1.330000 ;
      RECT 0.945000  2.185000 1.795000 2.635000 ;
      RECT 1.105000  1.330000 1.275000 1.785000 ;
      RECT 1.105000  1.785000 2.225000 2.005000 ;
      RECT 1.465000  0.255000 1.795000 0.635000 ;
      RECT 1.965000  0.465000 2.175000 0.635000 ;
      RECT 1.965000  0.635000 3.120000 0.825000 ;
      RECT 1.965000  2.005000 2.225000 2.465000 ;
      RECT 2.345000  0.085000 2.675000 0.465000 ;
      RECT 2.795000  1.650000 3.120000 2.635000 ;
      RECT 2.845000  0.495000 3.120000 0.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o21a_2
MACRO sky130_fd_sc_hd__o21a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.480000 0.990000 3.785000 1.495000 ;
        RECT 3.480000 1.495000 5.400000 1.705000 ;
        RECT 5.030000 0.995000 5.400000 1.495000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.140000 0.995000 4.690000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485000 1.075000 3.155000 1.615000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.635000 1.715000 0.805000 ;
        RECT 0.090000 0.805000 0.320000 1.530000 ;
        RECT 0.090000 1.530000 1.955000 1.700000 ;
        RECT 0.595000 0.615000 1.715000 0.635000 ;
        RECT 0.915000 1.700000 1.105000 2.465000 ;
        RECT 1.775000 1.700000 1.955000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.415000  1.870000 0.745000 2.635000 ;
      RECT 0.490000  0.995000 2.315000 1.335000 ;
      RECT 0.955000  0.085000 1.285000 0.445000 ;
      RECT 1.275000  1.870000 1.605000 2.635000 ;
      RECT 1.815000  0.085000 2.145000 0.465000 ;
      RECT 2.115000  0.655000 3.095000 0.870000 ;
      RECT 2.115000  0.870000 2.315000 0.995000 ;
      RECT 2.125000  1.335000 2.315000 1.830000 ;
      RECT 2.125000  1.830000 2.845000 1.875000 ;
      RECT 2.125000  1.875000 4.545000 2.085000 ;
      RECT 2.135000  2.255000 2.485000 2.635000 ;
      RECT 2.335000  0.255000 3.605000 0.485000 ;
      RECT 2.655000  2.085000 4.545000 2.105000 ;
      RECT 2.655000  2.105000 2.845000 2.465000 ;
      RECT 3.015000  2.275000 3.685000 2.635000 ;
      RECT 3.275000  0.485000 3.605000 0.615000 ;
      RECT 3.275000  0.615000 5.405000 0.785000 ;
      RECT 3.775000  0.085000 4.115000 0.445000 ;
      RECT 4.215000  2.105000 4.545000 2.445000 ;
      RECT 4.645000  0.085000 4.975000 0.445000 ;
      RECT 5.075000  1.935000 5.435000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__o21a_4
MACRO sky130_fd_sc_hd__o21ai_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ai_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.415000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.100000 1.005000 1.340000 ;
        RECT 0.605000 1.340000 0.775000 1.645000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 1.355000 1.730000 1.685000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.290500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 1.510000 1.345000 1.680000 ;
        RECT 0.965000 1.680000 1.300000 2.465000 ;
        RECT 1.175000 0.955000 1.740000 1.125000 ;
        RECT 1.175000 1.125000 1.345000 1.510000 ;
        RECT 1.455000 0.280000 1.740000 0.955000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.120000  0.280000 0.380000 0.615000 ;
      RECT 0.120000  0.615000 1.285000 0.785000 ;
      RECT 0.145000  1.825000 0.475000 2.635000 ;
      RECT 0.550000  0.085000 0.880000 0.445000 ;
      RECT 1.050000  0.280000 1.285000 0.615000 ;
      RECT 1.470000  1.855000 1.725000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__o21ai_0
MACRO sky130_fd_sc_hd__o21ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.995000 0.410000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.590000 0.995000 0.975000 1.325000 ;
        RECT 0.590000 1.325000 0.785000 2.375000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.202500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.295000 1.750000 1.655000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.517000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 1.505000 1.315000 1.785000 ;
        RECT 0.965000 1.785000 1.295000 2.465000 ;
        RECT 1.145000 0.955000 1.665000 1.125000 ;
        RECT 1.145000 1.125000 1.315000 1.505000 ;
        RECT 1.495000 0.390000 1.665000 0.955000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.090000  0.265000 0.380000 0.615000 ;
      RECT 0.090000  0.615000 1.305000 0.785000 ;
      RECT 0.090000  1.495000 0.410000 2.635000 ;
      RECT 0.575000  0.085000 0.905000 0.445000 ;
      RECT 1.075000  0.310000 1.305000 0.615000 ;
      RECT 1.495000  1.835000 1.750000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__o21ai_1
MACRO sky130_fd_sc_hd__o21ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 1.055000 0.450000 1.445000 ;
        RECT 0.120000 1.445000 2.095000 1.615000 ;
        RECT 1.600000 1.075000 2.095000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.620000 1.075000 1.420000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.815000 0.765000 3.130000 1.400000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.742000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 1.785000 2.645000 1.965000 ;
        RECT 0.995000 1.965000 1.295000 2.125000 ;
        RECT 2.410000 1.965000 2.645000 2.465000 ;
        RECT 2.435000 0.595000 2.645000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.085000 0.310000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.105000  0.255000 0.435000 0.715000 ;
      RECT 0.105000  0.715000 2.265000 0.885000 ;
      RECT 0.105000  1.785000 0.435000 2.635000 ;
      RECT 0.605000  1.785000 0.825000 2.295000 ;
      RECT 0.605000  2.295000 1.715000 2.465000 ;
      RECT 0.615000  0.085000 0.785000 0.545000 ;
      RECT 0.965000  0.255000 1.295000 0.715000 ;
      RECT 1.525000  0.085000 1.695000 0.545000 ;
      RECT 1.525000  2.135000 1.715000 2.295000 ;
      RECT 1.910000  2.175000 2.240000 2.635000 ;
      RECT 1.935000  0.255000 3.125000 0.425000 ;
      RECT 1.935000  0.425000 2.265000 0.715000 ;
      RECT 2.815000  0.425000 3.125000 0.595000 ;
      RECT 2.815000  1.570000 3.125000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o21ai_2
MACRO sky130_fd_sc_hd__o21ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.015000 1.475000 1.320000 ;
        RECT 0.575000 1.320000 1.475000 1.515000 ;
        RECT 0.575000 1.515000 3.695000 1.685000 ;
        RECT 3.445000 0.990000 3.695000 1.515000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 1.070000 3.275000 1.345000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.905000 1.015000 5.255000 1.275000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.484000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.840000 1.855000 5.150000 2.025000 ;
        RECT 3.935000 1.445000 5.835000 1.700000 ;
        RECT 3.935000 1.700000 5.150000 1.855000 ;
        RECT 4.030000 0.615000 5.835000 0.845000 ;
        RECT 4.080000 2.025000 5.150000 2.085000 ;
        RECT 4.080000 2.085000 4.290000 2.465000 ;
        RECT 4.960000 2.085000 5.150000 2.465000 ;
        RECT 5.425000 0.845000 5.835000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.120000  0.615000 3.860000 0.820000 ;
      RECT 0.120000  1.820000 0.405000 2.635000 ;
      RECT 0.550000  0.085000 0.880000 0.445000 ;
      RECT 0.575000  1.915000 1.670000 2.085000 ;
      RECT 0.575000  2.085000 0.810000 2.465000 ;
      RECT 0.980000  2.255000 1.310000 2.635000 ;
      RECT 1.410000  0.085000 1.740000 0.445000 ;
      RECT 1.480000  2.085000 1.670000 2.275000 ;
      RECT 1.480000  2.275000 3.460000 2.465000 ;
      RECT 2.270000  0.085000 2.600000 0.445000 ;
      RECT 3.130000  0.085000 3.460000 0.445000 ;
      RECT 3.630000  0.255000 5.650000 0.445000 ;
      RECT 3.630000  0.445000 3.860000 0.615000 ;
      RECT 3.630000  2.195000 3.910000 2.635000 ;
      RECT 4.460000  2.255000 4.790000 2.635000 ;
      RECT 5.320000  1.880000 5.650000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__o21ai_4
MACRO sky130_fd_sc_hd__o21ba_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ba_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.950000 1.075000 3.595000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.210000 1.075000 2.780000 1.285000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.030000 0.995000 1.360000 1.325000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.450000 0.445000 0.825000 ;
        RECT 0.085000 0.825000 0.340000 1.480000 ;
        RECT 0.085000 1.480000 0.425000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.510000  0.995000 0.860000 1.325000 ;
      RECT 0.595000  1.325000 0.860000 1.865000 ;
      RECT 0.595000  1.865000 2.575000 2.035000 ;
      RECT 0.595000  2.205000 1.005000 2.635000 ;
      RECT 0.710000  0.085000 0.880000 0.825000 ;
      RECT 1.075000  1.525000 1.700000 1.695000 ;
      RECT 1.160000  0.450000 1.330000 0.655000 ;
      RECT 1.160000  0.655000 1.700000 0.825000 ;
      RECT 1.530000  0.825000 1.700000 1.525000 ;
      RECT 1.750000  2.215000 2.080000 2.635000 ;
      RECT 1.870000  0.255000 2.040000 1.455000 ;
      RECT 1.870000  1.455000 2.575000 1.865000 ;
      RECT 2.250000  2.035000 2.575000 2.465000 ;
      RECT 2.270000  0.255000 2.600000 0.735000 ;
      RECT 2.270000  0.735000 3.440000 0.905000 ;
      RECT 2.770000  0.085000 2.940000 0.555000 ;
      RECT 3.050000  1.535000 3.380000 2.635000 ;
      RECT 3.110000  0.270000 3.440000 0.735000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o21ba_1
MACRO sky130_fd_sc_hd__o21ba_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ba_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.100000 1.075000 3.595000 1.625000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.075000 2.930000 1.285000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.325000 ;
        RECT 0.595000 1.325000 0.775000 1.695000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.255000 1.240000 0.595000 ;
        RECT 0.945000 0.595000 1.115000 1.495000 ;
        RECT 0.945000 1.495000 1.350000 1.695000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.430000 0.345000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.495000 ;
      RECT 0.085000  1.495000 0.395000 1.865000 ;
      RECT 0.085000  1.865000 1.935000 2.035000 ;
      RECT 0.520000  2.205000 0.910000 2.635000 ;
      RECT 0.595000  0.085000 0.775000 0.825000 ;
      RECT 1.285000  0.890000 1.595000 1.060000 ;
      RECT 1.285000  1.060000 1.455000 1.325000 ;
      RECT 1.410000  0.085000 1.770000 0.485000 ;
      RECT 1.415000  2.205000 2.230000 2.635000 ;
      RECT 1.425000  0.655000 2.275000 0.825000 ;
      RECT 1.425000  0.825000 1.595000 0.890000 ;
      RECT 1.765000  0.995000 1.935000 1.865000 ;
      RECT 1.940000  0.255000 2.275000 0.655000 ;
      RECT 2.105000  0.825000 2.275000 1.455000 ;
      RECT 2.105000  1.455000 2.725000 2.035000 ;
      RECT 2.400000  2.035000 2.725000 2.465000 ;
      RECT 2.445000  0.365000 2.745000 0.735000 ;
      RECT 2.445000  0.735000 3.590000 0.905000 ;
      RECT 2.915000  0.085000 3.085000 0.555000 ;
      RECT 3.200000  1.875000 3.530000 2.635000 ;
      RECT 3.255000  0.270000 3.590000 0.735000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o21ba_2
MACRO sky130_fd_sc_hd__o21ba_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ba_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.990000 1.075000 5.895000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.780000 1.075000 4.820000 1.275000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 0.885000 1.285000 ;
        RECT 0.605000 1.285000 0.885000 1.705000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 0.255000 1.385000 0.725000 ;
        RECT 1.055000 0.725000 2.225000 0.905000 ;
        RECT 1.055000 0.905000 1.455000 1.445000 ;
        RECT 1.055000 1.445000 2.225000 1.705000 ;
        RECT 1.895000 0.255000 2.225000 0.725000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.265000 0.545000 0.855000 ;
      RECT 0.085000  0.855000 0.255000 1.455000 ;
      RECT 0.085000  1.455000 0.435000 1.875000 ;
      RECT 0.085000  1.875000 2.565000 2.045000 ;
      RECT 0.085000  2.045000 0.435000 2.465000 ;
      RECT 0.635000  2.215000 0.965000 2.635000 ;
      RECT 0.715000  0.085000 0.885000 0.905000 ;
      RECT 1.475000  2.215000 1.805000 2.635000 ;
      RECT 1.555000  0.085000 1.725000 0.555000 ;
      RECT 1.625000  1.075000 2.565000 1.275000 ;
      RECT 2.315000  2.215000 2.645000 2.635000 ;
      RECT 2.395000  0.085000 2.565000 0.555000 ;
      RECT 2.395000  0.725000 3.585000 0.895000 ;
      RECT 2.395000  0.895000 2.565000 1.075000 ;
      RECT 2.395000  1.445000 2.905000 1.615000 ;
      RECT 2.395000  1.615000 2.565000 1.875000 ;
      RECT 2.735000  1.075000 3.135000 1.245000 ;
      RECT 2.735000  1.245000 2.905000 1.445000 ;
      RECT 2.805000  0.255000 4.005000 0.475000 ;
      RECT 2.815000  1.795000 4.380000 1.965000 ;
      RECT 2.815000  1.965000 2.985000 2.465000 ;
      RECT 3.200000  2.135000 3.450000 2.635000 ;
      RECT 3.235000  0.645000 3.585000 0.725000 ;
      RECT 3.395000  0.895000 3.585000 1.795000 ;
      RECT 3.685000  2.135000 3.925000 2.295000 ;
      RECT 3.685000  2.295000 4.765000 2.465000 ;
      RECT 3.755000  0.475000 4.005000 0.725000 ;
      RECT 3.755000  0.725000 5.710000 0.905000 ;
      RECT 4.135000  1.445000 4.380000 1.795000 ;
      RECT 4.135000  1.965000 4.380000 2.125000 ;
      RECT 4.175000  0.085000 4.345000 0.555000 ;
      RECT 4.515000  0.255000 4.845000 0.725000 ;
      RECT 4.595000  1.455000 5.710000 1.665000 ;
      RECT 4.595000  1.665000 4.765000 2.295000 ;
      RECT 4.935000  1.835000 5.265000 2.635000 ;
      RECT 5.015000  0.085000 5.185000 0.555000 ;
      RECT 5.355000  0.265000 5.710000 0.725000 ;
      RECT 5.435000  1.665000 5.710000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__o21ba_4
MACRO sky130_fd_sc_hd__o21bai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21bai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195000 1.075000 2.675000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 1.075000 2.025000 1.285000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.535000 1.345000 ;
        RECT 0.085000 1.345000 0.355000 2.445000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.474000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 0.255000 1.285000 0.645000 ;
        RECT 1.115000 0.645000 1.355000 0.825000 ;
        RECT 1.185000 0.825000 1.355000 1.455000 ;
        RECT 1.185000 1.455000 1.795000 1.625000 ;
        RECT 1.470000 1.625000 1.795000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.085000 0.360000 0.825000 ;
      RECT 0.525000  1.535000 1.015000 1.705000 ;
      RECT 0.525000  1.705000 0.800000 2.210000 ;
      RECT 0.580000  0.495000 0.770000 0.655000 ;
      RECT 0.580000  0.655000 0.890000 0.825000 ;
      RECT 0.720000  0.825000 0.890000 0.995000 ;
      RECT 0.720000  0.995000 1.015000 1.535000 ;
      RECT 0.970000  1.875000 1.300000 2.635000 ;
      RECT 1.490000  0.255000 1.820000 0.485000 ;
      RECT 1.570000  0.485000 1.740000 0.735000 ;
      RECT 1.570000  0.735000 2.665000 0.905000 ;
      RECT 1.995000  0.085000 2.165000 0.555000 ;
      RECT 2.270000  1.535000 2.645000 2.635000 ;
      RECT 2.335000  0.270000 2.665000 0.735000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__o21bai_1
MACRO sky130_fd_sc_hd__o21bai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21bai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.260000 1.075000 4.055000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.950000 1.075000 3.090000 1.275000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.525000 1.325000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.445000 2.650000 1.615000 ;
        RECT 1.085000 1.615000 1.255000 2.465000 ;
        RECT 1.525000 0.645000 1.855000 0.905000 ;
        RECT 1.525000 0.905000 1.780000 1.445000 ;
        RECT 2.405000 1.615000 2.650000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.180000  0.085000 0.350000 0.825000 ;
      RECT 0.180000  1.495000 0.865000 1.665000 ;
      RECT 0.180000  1.665000 0.350000 1.915000 ;
      RECT 0.585000  1.875000 0.915000 2.635000 ;
      RECT 0.600000  0.445000 0.865000 0.825000 ;
      RECT 0.695000  0.825000 0.865000 1.075000 ;
      RECT 0.695000  1.075000 1.335000 1.245000 ;
      RECT 0.695000  1.245000 0.865000 1.495000 ;
      RECT 1.075000  0.255000 2.275000 0.475000 ;
      RECT 1.075000  0.475000 1.355000 0.905000 ;
      RECT 1.470000  1.795000 1.720000 2.635000 ;
      RECT 1.955000  1.795000 2.235000 2.295000 ;
      RECT 1.955000  2.295000 3.035000 2.465000 ;
      RECT 2.025000  0.475000 2.275000 0.725000 ;
      RECT 2.025000  0.725000 3.980000 0.905000 ;
      RECT 2.445000  0.085000 2.615000 0.555000 ;
      RECT 2.785000  0.255000 3.115000 0.725000 ;
      RECT 2.865000  1.455000 3.980000 1.665000 ;
      RECT 2.865000  1.665000 3.035000 2.295000 ;
      RECT 3.205000  1.835000 3.535000 2.635000 ;
      RECT 3.285000  0.085000 3.455000 0.555000 ;
      RECT 3.625000  0.265000 3.980000 0.725000 ;
      RECT 3.705000  1.665000 3.980000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__o21bai_2
MACRO sky130_fd_sc_hd__o21bai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21bai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.645000 1.075000 6.810000 1.285000 ;
        RECT 6.585000 1.285000 6.810000 2.455000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.065000 1.075000 4.475000 1.275000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.555000 1.285000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.455000 4.315000 1.625000 ;
        RECT 1.065000 1.625000 1.275000 2.465000 ;
        RECT 1.420000 0.645000 2.675000 0.815000 ;
        RECT 1.865000 1.625000 2.115000 2.465000 ;
        RECT 2.445000 0.815000 2.675000 1.075000 ;
        RECT 2.445000 1.075000 2.895000 1.445000 ;
        RECT 2.445000 1.445000 4.315000 1.455000 ;
        RECT 3.225000 1.625000 3.475000 2.125000 ;
        RECT 4.065000 1.625000 4.315000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.090000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.145000  1.455000 0.895000 1.625000 ;
      RECT 0.145000  1.625000 0.475000 2.435000 ;
      RECT 0.225000  0.085000 0.395000 0.895000 ;
      RECT 0.565000  0.290000 0.895000 0.895000 ;
      RECT 0.645000  1.795000 0.855000 2.635000 ;
      RECT 0.725000  0.895000 0.895000 1.075000 ;
      RECT 0.725000  1.075000 2.275000 1.285000 ;
      RECT 0.725000  1.285000 0.895000 1.455000 ;
      RECT 1.080000  0.305000 3.095000 0.475000 ;
      RECT 1.445000  1.795000 1.695000 2.635000 ;
      RECT 2.285000  1.795000 2.535000 2.635000 ;
      RECT 2.775000  1.795000 3.055000 2.295000 ;
      RECT 2.775000  2.295000 4.735000 2.465000 ;
      RECT 2.845000  0.475000 3.095000 0.725000 ;
      RECT 2.845000  0.725000 6.455000 0.905000 ;
      RECT 3.265000  0.085000 3.435000 0.555000 ;
      RECT 3.605000  0.255000 3.935000 0.725000 ;
      RECT 3.645000  1.795000 3.895000 2.295000 ;
      RECT 4.105000  0.085000 4.275000 0.555000 ;
      RECT 4.445000  0.255000 4.775000 0.725000 ;
      RECT 4.485000  1.455000 6.415000 1.625000 ;
      RECT 4.485000  1.625000 4.735000 2.295000 ;
      RECT 4.905000  1.795000 5.155000 2.635000 ;
      RECT 4.945000  0.085000 5.115000 0.555000 ;
      RECT 5.285000  0.255000 5.615000 0.725000 ;
      RECT 5.325000  1.625000 5.575000 2.465000 ;
      RECT 5.745000  1.795000 5.995000 2.635000 ;
      RECT 5.785000  0.085000 5.955000 0.555000 ;
      RECT 6.125000  0.255000 6.455000 0.725000 ;
      RECT 6.165000  1.625000 6.415000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
END sky130_fd_sc_hd__o21bai_4
MACRO sky130_fd_sc_hd__o22a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.670000 1.075000 3.135000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.165000 1.075000 2.495000 1.325000 ;
        RECT 2.315000 1.325000 2.495000 1.445000 ;
        RECT 2.315000 1.445000 2.645000 1.615000 ;
        RECT 2.445000 1.615000 2.645000 2.405000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.980000 1.075000 1.335000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 1.075000 1.995000 1.325000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.365000 0.365000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.535000  0.715000 1.785000 0.895000 ;
      RECT 0.535000  0.895000 0.810000 1.495000 ;
      RECT 0.535000  1.495000 2.145000 1.705000 ;
      RECT 0.555000  1.875000 1.340000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.545000 ;
      RECT 1.035000  0.295000 2.285000 0.475000 ;
      RECT 1.420000  0.645000 1.785000 0.715000 ;
      RECT 1.735000  1.705000 2.145000 1.805000 ;
      RECT 1.735000  1.805000 2.120000 2.465000 ;
      RECT 1.955000  0.475000 2.285000 0.695000 ;
      RECT 1.955000  0.695000 3.135000 0.865000 ;
      RECT 2.455000  0.085000 2.625000 0.525000 ;
      RECT 2.795000  0.280000 3.135000 0.695000 ;
      RECT 2.815000  1.455000 3.135000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o22a_1
MACRO sky130_fd_sc_hd__o22a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095000 1.075000 3.590000 1.275000 ;
        RECT 3.270000 1.275000 3.590000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.595000 1.075000 2.925000 1.325000 ;
        RECT 2.745000 1.325000 2.925000 1.445000 ;
        RECT 2.745000 1.445000 3.100000 1.615000 ;
        RECT 2.900000 1.615000 3.100000 2.405000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 1.075000 1.790000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.960000 1.075000 2.425000 1.325000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.590000 0.365000 0.805000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.130000 -0.085000 0.300000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.115000  1.445000 0.365000 2.635000 ;
      RECT 0.185000  0.085000 0.355000 0.885000 ;
      RECT 0.975000  0.715000 2.215000 0.895000 ;
      RECT 0.975000  0.895000 1.255000 1.495000 ;
      RECT 0.975000  1.495000 2.575000 1.705000 ;
      RECT 0.995000  1.875000 1.795000 2.635000 ;
      RECT 1.025000  0.085000 1.205000 0.545000 ;
      RECT 1.465000  0.295000 2.730000 0.475000 ;
      RECT 1.850000  0.645000 2.215000 0.715000 ;
      RECT 2.190000  1.705000 2.575000 2.465000 ;
      RECT 2.390000  0.475000 2.730000 0.695000 ;
      RECT 2.390000  0.695000 3.590000 0.825000 ;
      RECT 2.560000  0.825000 3.590000 0.865000 ;
      RECT 2.915000  0.085000 3.085000 0.525000 ;
      RECT 3.255000  0.280000 3.590000 0.695000 ;
      RECT 3.270000  1.795000 3.590000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o22a_2
MACRO sky130_fd_sc_hd__o22a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.350000 1.075000 4.680000 1.445000 ;
        RECT 4.350000 1.445000 5.735000 1.615000 ;
        RECT 5.565000 1.075000 6.355000 1.275000 ;
        RECT 5.565000 1.275000 5.735000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.900000 1.075000 5.395000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.420000 1.075000 2.955000 1.445000 ;
        RECT 2.420000 1.445000 4.180000 1.615000 ;
        RECT 3.850000 1.075000 4.180000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.125000 1.075000 3.680000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.725000 1.770000 0.905000 ;
        RECT 0.085000 0.905000 0.370000 1.445000 ;
        RECT 0.085000 1.445000 1.730000 1.615000 ;
        RECT 0.600000 0.265000 0.930000 0.725000 ;
        RECT 0.640000 1.615000 0.890000 2.465000 ;
        RECT 1.440000 0.255000 1.770000 0.725000 ;
        RECT 1.480000 1.615000 1.730000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.220000  1.825000 0.470000 2.635000 ;
      RECT 0.260000  0.085000 0.430000 0.555000 ;
      RECT 0.540000  1.075000 2.230000 1.275000 ;
      RECT 1.060000  1.795000 1.310000 2.635000 ;
      RECT 1.100000  0.085000 1.270000 0.555000 ;
      RECT 1.900000  1.275000 2.230000 1.785000 ;
      RECT 1.900000  1.785000 5.270000 1.955000 ;
      RECT 1.900000  2.125000 2.670000 2.635000 ;
      RECT 1.940000  0.085000 2.110000 0.555000 ;
      RECT 1.940000  0.735000 3.970000 0.905000 ;
      RECT 1.940000  0.905000 2.230000 1.075000 ;
      RECT 2.380000  0.255000 4.470000 0.475000 ;
      RECT 2.415000  0.645000 3.970000 0.735000 ;
      RECT 2.840000  2.125000 3.090000 2.295000 ;
      RECT 2.840000  2.295000 3.930000 2.465000 ;
      RECT 3.260000  1.955000 3.510000 2.125000 ;
      RECT 3.680000  2.125000 3.930000 2.295000 ;
      RECT 4.100000  2.125000 4.430000 2.635000 ;
      RECT 4.140000  0.475000 4.470000 0.735000 ;
      RECT 4.140000  0.735000 6.150000 0.905000 ;
      RECT 4.600000  2.125000 4.850000 2.295000 ;
      RECT 4.600000  2.295000 5.690000 2.465000 ;
      RECT 4.640000  0.085000 4.810000 0.555000 ;
      RECT 4.980000  0.255000 5.310000 0.725000 ;
      RECT 4.980000  0.725000 6.150000 0.735000 ;
      RECT 5.020000  1.955000 5.270000 2.125000 ;
      RECT 5.440000  1.785000 5.690000 2.295000 ;
      RECT 5.480000  0.085000 5.650000 0.555000 ;
      RECT 5.820000  0.255000 6.150000 0.725000 ;
      RECT 5.905000  1.455000 6.110000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__o22a_4
MACRO sky130_fd_sc_hd__o22ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.755000 1.075000 2.215000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.220000 1.075000 1.585000 1.245000 ;
        RECT 1.405000 1.245000 1.585000 1.445000 ;
        RECT 1.405000 1.445000 1.725000 1.615000 ;
        RECT 1.525000 1.615000 1.725000 2.405000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.665000 0.325000 1.990000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835000 0.995000 1.005000 1.415000 ;
        RECT 0.835000 1.415000 1.235000 1.665000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.650250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.495000 0.645000 0.845000 0.825000 ;
        RECT 0.495000 0.825000 0.665000 1.835000 ;
        RECT 0.495000 1.835000 1.335000 2.045000 ;
        RECT 0.835000 2.045000 1.335000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.085000  0.295000 1.345000 0.475000 ;
      RECT 0.135000  2.175000 0.345000 2.635000 ;
      RECT 1.015000  0.475000 1.345000 0.695000 ;
      RECT 1.015000  0.695000 2.215000 0.825000 ;
      RECT 1.185000  0.825000 2.215000 0.865000 ;
      RECT 1.535000  0.085000 1.705000 0.525000 ;
      RECT 1.875000  0.280000 2.215000 0.695000 ;
      RECT 1.895000  1.455000 2.215000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__o22ai_1
MACRO sky130_fd_sc_hd__o22ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395000 1.075000 4.165000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.075000 3.225000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.200000 1.075000 0.985000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.155000 1.075000 1.925000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.645000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 2.340000 0.905000 ;
        RECT 1.375000 0.645000 1.705000 0.725000 ;
        RECT 1.415000 1.445000 3.065000 1.625000 ;
        RECT 1.415000 1.625000 1.665000 2.125000 ;
        RECT 2.095000 0.905000 2.340000 1.445000 ;
        RECT 2.815000 1.625000 3.065000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  0.305000 2.680000 0.475000 ;
      RECT 0.090000  0.475000 0.365000 0.905000 ;
      RECT 0.150000  1.455000 1.245000 1.625000 ;
      RECT 0.150000  1.625000 0.405000 2.465000 ;
      RECT 0.575000  1.795000 0.825000 2.635000 ;
      RECT 0.995000  1.625000 1.245000 2.295000 ;
      RECT 0.995000  2.295000 2.085000 2.465000 ;
      RECT 1.835000  1.795000 2.085000 2.295000 ;
      RECT 2.395000  1.795000 2.645000 2.295000 ;
      RECT 2.395000  2.295000 3.485000 2.465000 ;
      RECT 2.510000  0.475000 2.680000 0.725000 ;
      RECT 2.510000  0.725000 4.365000 0.905000 ;
      RECT 2.855000  0.085000 3.025000 0.555000 ;
      RECT 3.195000  0.255000 3.525000 0.725000 ;
      RECT 3.235000  1.455000 4.330000 1.625000 ;
      RECT 3.235000  1.625000 3.485000 2.295000 ;
      RECT 3.655000  1.795000 3.905000 2.635000 ;
      RECT 3.695000  0.085000 3.865000 0.555000 ;
      RECT 4.035000  0.255000 4.365000 0.725000 ;
      RECT 4.075000  1.625000 4.330000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__o22ai_2
MACRO sky130_fd_sc_hd__o22ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 1.415000 1.275000 ;
        RECT 1.150000 1.275000 1.415000 1.445000 ;
        RECT 1.150000 1.445000 3.575000 1.615000 ;
        RECT 3.275000 1.075000 3.605000 1.245000 ;
        RECT 3.275000 1.245000 3.575000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.685000 1.075000 3.095000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.295000 0.995000 4.940000 1.445000 ;
        RECT 4.295000 1.445000 6.935000 1.615000 ;
        RECT 6.715000 0.995000 6.935000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.110000 1.075000 6.460000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.845000 1.785000 3.915000 1.955000 ;
        RECT 1.845000 1.955000 2.095000 2.125000 ;
        RECT 2.685000 1.955000 2.935000 2.125000 ;
        RECT 3.745000 1.445000 4.125000 1.615000 ;
        RECT 3.745000 1.615000 3.915000 1.785000 ;
        RECT 3.955000 0.645000 7.275000 0.820000 ;
        RECT 3.955000 0.820000 4.125000 1.445000 ;
        RECT 5.255000 1.785000 7.275000 1.955000 ;
        RECT 5.255000 1.955000 5.505000 2.125000 ;
        RECT 6.095000 1.955000 6.345000 2.125000 ;
        RECT 7.105000 0.820000 7.275000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.125000  0.255000 0.455000 0.725000 ;
      RECT 0.125000  0.725000 1.295000 0.735000 ;
      RECT 0.125000  0.735000 3.785000 0.905000 ;
      RECT 0.165000  1.445000 0.415000 2.635000 ;
      RECT 0.585000  1.445000 0.835000 1.785000 ;
      RECT 0.585000  1.785000 1.675000 1.955000 ;
      RECT 0.585000  1.955000 0.835000 2.465000 ;
      RECT 0.625000  0.085000 0.795000 0.555000 ;
      RECT 0.965000  0.255000 1.295000 0.725000 ;
      RECT 1.005000  2.125000 1.255000 2.635000 ;
      RECT 1.425000  1.955000 1.675000 2.295000 ;
      RECT 1.425000  2.295000 3.395000 2.465000 ;
      RECT 1.465000  0.085000 1.635000 0.555000 ;
      RECT 1.805000  0.255000 2.135000 0.725000 ;
      RECT 1.805000  0.725000 2.975000 0.735000 ;
      RECT 2.265000  2.125000 2.515000 2.295000 ;
      RECT 2.305000  0.085000 2.475000 0.555000 ;
      RECT 2.645000  0.255000 2.975000 0.725000 ;
      RECT 3.105000  2.125000 3.395000 2.295000 ;
      RECT 3.145000  0.085000 3.315000 0.555000 ;
      RECT 3.485000  0.255000 7.245000 0.475000 ;
      RECT 3.485000  0.475000 3.785000 0.735000 ;
      RECT 3.565000  2.125000 3.785000 2.635000 ;
      RECT 3.955000  2.125000 4.255000 2.465000 ;
      RECT 4.085000  1.785000 5.085000 1.955000 ;
      RECT 4.085000  1.955000 4.255000 2.125000 ;
      RECT 4.425000  2.125000 4.665000 2.635000 ;
      RECT 4.835000  1.955000 5.085000 2.295000 ;
      RECT 4.835000  2.295000 6.765000 2.465000 ;
      RECT 5.675000  2.125000 5.925000 2.295000 ;
      RECT 6.515000  2.135000 6.765000 2.295000 ;
      RECT 6.935000  2.125000 7.215000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__o22ai_4
MACRO sky130_fd_sc_hd__o31a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.905000 0.995000 1.295000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 0.995000 1.725000 1.325000 ;
        RECT 1.525000 1.325000 1.725000 2.125000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925000 0.995000 2.175000 2.125000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.390000 0.995000 2.795000 1.325000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.594000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.265000 0.525000 0.825000 ;
        RECT 0.085000 0.825000 0.395000 1.835000 ;
        RECT 0.085000 1.835000 0.525000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.565000  0.995000 0.735000 1.445000 ;
      RECT 0.565000  1.445000 1.355000 1.615000 ;
      RECT 0.695000  0.085000 1.145000 0.825000 ;
      RECT 0.700000  1.785000 1.015000 2.635000 ;
      RECT 1.185000  1.615000 1.355000 2.295000 ;
      RECT 1.185000  2.295000 2.615000 2.465000 ;
      RECT 1.315000  0.255000 1.485000 0.655000 ;
      RECT 1.315000  0.655000 2.475000 0.825000 ;
      RECT 1.655000  0.085000 2.075000 0.485000 ;
      RECT 2.245000  0.255000 2.475000 0.655000 ;
      RECT 2.365000  1.495000 3.135000 1.665000 ;
      RECT 2.365000  1.665000 2.615000 2.295000 ;
      RECT 2.645000  0.255000 3.135000 0.825000 ;
      RECT 2.795000  1.835000 3.125000 2.635000 ;
      RECT 2.965000  0.825000 3.135000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o31a_1
MACRO sky130_fd_sc_hd__o31a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.370000 0.995000 1.760000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 0.995000 2.190000 1.325000 ;
        RECT 1.990000 1.325000 2.190000 2.125000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.390000 0.995000 2.640000 2.125000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855000 0.995000 3.255000 1.325000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.577500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.860000 1.295000 ;
        RECT 0.550000 0.265000 0.990000 0.825000 ;
        RECT 0.550000 0.825000 0.860000 1.075000 ;
        RECT 0.550000 1.295000 0.860000 1.835000 ;
        RECT 0.550000 1.835000 0.990000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.085000 0.380000 0.905000 ;
      RECT 0.085000  1.465000 0.380000 2.635000 ;
      RECT 1.030000  0.995000 1.200000 1.445000 ;
      RECT 1.030000  1.445000 1.820000 1.615000 ;
      RECT 1.160000  0.085000 1.610000 0.825000 ;
      RECT 1.165000  1.785000 1.480000 2.635000 ;
      RECT 1.650000  1.615000 1.820000 2.295000 ;
      RECT 1.650000  2.295000 3.080000 2.465000 ;
      RECT 1.780000  0.255000 1.950000 0.655000 ;
      RECT 1.780000  0.655000 2.940000 0.825000 ;
      RECT 2.120000  0.085000 2.540000 0.485000 ;
      RECT 2.710000  0.255000 2.940000 0.655000 ;
      RECT 2.830000  1.495000 3.595000 1.665000 ;
      RECT 2.830000  1.665000 3.080000 2.295000 ;
      RECT 3.110000  0.255000 3.595000 0.825000 ;
      RECT 3.255000  1.835000 3.590000 2.635000 ;
      RECT 3.425000  0.825000 3.595000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o31a_2
MACRO sky130_fd_sc_hd__o31a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.140000 1.055000 5.470000 1.360000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.265000 1.055000 4.970000 1.360000 ;
        RECT 4.680000 1.360000 4.970000 1.530000 ;
        RECT 4.680000 1.530000 6.355000 1.700000 ;
        RECT 5.640000 1.055000 6.355000 1.530000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765000 1.055000 4.095000 1.360000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.780000 1.055000 3.575000 1.355000 ;
        RECT 2.780000 1.355000 3.150000 1.695000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 1.765000 0.885000 ;
        RECT 0.085000 0.885000 0.735000 1.460000 ;
        RECT 0.085000 1.460000 1.750000 1.665000 ;
        RECT 0.680000 0.255000 0.895000 0.655000 ;
        RECT 0.680000 0.655000 1.765000 0.715000 ;
        RECT 0.680000 1.665000 0.895000 2.465000 ;
        RECT 1.565000 0.255000 1.765000 0.655000 ;
        RECT 1.565000 1.665000 1.750000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.125000 -0.085000 0.295000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.085000  0.085000 0.510000 0.545000 ;
      RECT 0.085000  1.835000 0.510000 2.635000 ;
      RECT 0.905000  1.055000 2.610000 1.290000 ;
      RECT 1.065000  0.085000 1.395000 0.485000 ;
      RECT 1.065000  1.835000 1.395000 2.635000 ;
      RECT 1.920000  1.460000 2.250000 2.635000 ;
      RECT 1.935000  0.085000 2.250000 0.885000 ;
      RECT 2.440000  0.255000 3.570000 0.465000 ;
      RECT 2.440000  0.635000 3.210000 0.885000 ;
      RECT 2.440000  0.885000 2.610000 1.055000 ;
      RECT 2.440000  1.290000 2.610000 1.870000 ;
      RECT 2.440000  1.870000 4.090000 2.070000 ;
      RECT 2.440000  2.070000 2.610000 2.465000 ;
      RECT 2.780000  2.240000 3.110000 2.635000 ;
      RECT 3.320000  1.530000 4.510000 1.700000 ;
      RECT 3.380000  0.465000 3.570000 0.635000 ;
      RECT 3.380000  0.635000 6.355000 0.885000 ;
      RECT 3.760000  0.085000 4.090000 0.445000 ;
      RECT 3.760000  2.070000 4.090000 2.465000 ;
      RECT 4.260000  0.255000 4.430000 0.635000 ;
      RECT 4.260000  1.700000 4.510000 2.465000 ;
      RECT 4.600000  0.085000 4.930000 0.445000 ;
      RECT 4.680000  1.870000 5.720000 2.070000 ;
      RECT 4.680000  2.070000 4.850000 2.465000 ;
      RECT 5.020000  2.240000 5.350000 2.635000 ;
      RECT 5.100000  0.255000 5.270000 0.635000 ;
      RECT 5.440000  0.085000 5.770000 0.445000 ;
      RECT 5.520000  2.070000 5.720000 2.465000 ;
      RECT 5.890000  1.870000 6.355000 2.465000 ;
      RECT 5.940000  0.255000 6.355000 0.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.125000 4.455000 2.295000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.125000 6.295000 2.295000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 4.225000 2.095000 4.515000 2.140000 ;
      RECT 4.225000 2.140000 6.355000 2.280000 ;
      RECT 4.225000 2.280000 4.515000 2.325000 ;
      RECT 6.065000 2.095000 6.355000 2.140000 ;
      RECT 6.065000 2.280000 6.355000 2.325000 ;
  END
END sky130_fd_sc_hd__o31a_4
MACRO sky130_fd_sc_hd__o31ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.440000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 1.075000 1.055000 2.465000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225000 1.075000 1.700000 1.325000 ;
        RECT 1.460000 1.325000 1.700000 2.405000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.330000 0.995000 2.675000 1.325000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.006000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 0.260000 2.675000 0.825000 ;
        RECT 1.945000 0.825000 2.160000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.090000  1.495000 0.440000 2.635000 ;
      RECT 0.175000  0.085000 0.345000 0.905000 ;
      RECT 0.515000  0.255000 0.845000 0.735000 ;
      RECT 0.515000  0.735000 1.700000 0.905000 ;
      RECT 1.015000  0.085000 1.185000 0.565000 ;
      RECT 1.370000  0.255000 1.700000 0.735000 ;
      RECT 2.330000  1.495000 2.675000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__o31ai_1
MACRO sky130_fd_sc_hd__o31ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.055000 1.240000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.410000 1.055000 2.220000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.390000 1.055000 3.205000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175000 0.755000 4.515000 1.325000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.063500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335000 1.495000 4.515000 1.665000 ;
        RECT 2.335000 1.665000 2.665000 2.125000 ;
        RECT 3.175000 1.665000 3.505000 2.465000 ;
        RECT 3.675000 0.595000 4.005000 1.495000 ;
        RECT 4.175000 1.665000 4.515000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  0.255000 0.445000 0.715000 ;
      RECT 0.090000  0.715000 3.505000 0.885000 ;
      RECT 0.090000  1.495000 2.125000 1.665000 ;
      RECT 0.090000  1.665000 0.445000 2.465000 ;
      RECT 0.615000  0.085000 0.785000 0.545000 ;
      RECT 0.615000  1.835000 0.785000 2.635000 ;
      RECT 0.955000  0.255000 1.285000 0.715000 ;
      RECT 0.955000  1.665000 1.285000 2.465000 ;
      RECT 1.455000  0.085000 1.965000 0.545000 ;
      RECT 1.455000  1.835000 1.625000 2.295000 ;
      RECT 1.455000  2.295000 3.005000 2.465000 ;
      RECT 1.795000  1.665000 2.125000 2.125000 ;
      RECT 2.175000  0.255000 2.505000 0.715000 ;
      RECT 2.675000  0.085000 3.005000 0.545000 ;
      RECT 2.835000  1.835000 3.005000 2.295000 ;
      RECT 3.175000  0.255000 4.515000 0.425000 ;
      RECT 3.175000  0.425000 3.505000 0.715000 ;
      RECT 3.675000  1.835000 4.005000 2.635000 ;
      RECT 4.175000  0.425000 4.515000 0.585000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__o31ai_2
MACRO sky130_fd_sc_hd__o31ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.055000 1.780000 1.425000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.950000 1.055000 3.605000 1.425000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775000 1.055000 5.940000 1.275000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.465000 1.055000 7.735000 1.275000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.683800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775000 1.445000 7.735000 1.695000 ;
        RECT 5.770000 1.695000 5.940000 2.465000 ;
        RECT 6.110000 0.645000 7.280000 0.885000 ;
        RECT 6.110000 0.885000 6.295000 1.445000 ;
        RECT 6.610000 1.695000 6.780000 2.465000 ;
        RECT 7.450000 1.695000 7.735000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.090000  0.255000 0.445000 0.715000 ;
      RECT 0.090000  0.715000 5.940000 0.885000 ;
      RECT 0.090000  1.595000 2.125000 1.895000 ;
      RECT 0.090000  1.895000 0.445000 2.465000 ;
      RECT 0.615000  0.085000 0.785000 0.545000 ;
      RECT 0.615000  2.065000 0.785000 2.635000 ;
      RECT 0.955000  0.255000 1.285000 0.715000 ;
      RECT 0.955000  1.895000 1.285000 2.465000 ;
      RECT 1.455000  0.085000 1.625000 0.545000 ;
      RECT 1.455000  2.065000 1.625000 2.635000 ;
      RECT 1.795000  0.255000 2.125000 0.715000 ;
      RECT 1.795000  1.895000 2.125000 2.205000 ;
      RECT 1.795000  2.205000 3.885000 2.465000 ;
      RECT 2.295000  0.085000 2.465000 0.545000 ;
      RECT 2.295000  1.595000 3.605000 1.765000 ;
      RECT 2.295000  1.765000 2.465000 2.035000 ;
      RECT 2.635000  0.255000 2.965000 0.715000 ;
      RECT 2.635000  1.935000 2.965000 2.205000 ;
      RECT 3.135000  0.085000 3.305000 0.545000 ;
      RECT 3.135000  1.765000 3.605000 1.865000 ;
      RECT 3.135000  1.865000 5.600000 2.035000 ;
      RECT 3.475000  0.255000 3.805000 0.715000 ;
      RECT 3.995000  0.085000 4.640000 0.545000 ;
      RECT 4.080000  2.035000 5.600000 2.465000 ;
      RECT 4.810000  0.395000 4.980000 0.715000 ;
      RECT 5.150000  0.085000 5.600000 0.545000 ;
      RECT 5.770000  0.255000 7.735000 0.475000 ;
      RECT 5.770000  0.475000 5.940000 0.715000 ;
      RECT 6.110000  1.890000 6.440000 2.635000 ;
      RECT 6.950000  1.890000 7.280000 2.635000 ;
      RECT 7.450000  0.475000 7.735000 0.885000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__o31ai_4
MACRO sky130_fd_sc_hd__o32a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 0.995000 1.175000 1.075000 ;
        RECT 1.005000 1.075000 1.255000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 0.995000 1.810000 1.325000 ;
        RECT 1.485000 1.325000 1.810000 2.125000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.980000 0.995000 2.255000 1.660000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.320000 0.995000 3.595000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.440000 0.995000 2.795000 1.660000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.504000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.595000 0.825000 ;
        RECT 0.085000 0.825000 0.260000 1.495000 ;
        RECT 0.085000 1.495000 0.470000 2.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.085000 0.310000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.445000  0.995000 0.635000 1.075000 ;
      RECT 0.445000  1.075000 0.810000 1.325000 ;
      RECT 0.640000  1.325000 0.810000 1.495000 ;
      RECT 0.640000  1.495000 1.315000 1.665000 ;
      RECT 0.685000  1.835000 0.975000 2.635000 ;
      RECT 0.765000  0.085000 0.935000 0.645000 ;
      RECT 1.140000  0.255000 1.470000 0.655000 ;
      RECT 1.140000  0.655000 2.540000 0.825000 ;
      RECT 1.145000  1.665000 1.315000 2.295000 ;
      RECT 1.145000  2.295000 2.510000 2.465000 ;
      RECT 1.645000  0.085000 1.975000 0.485000 ;
      RECT 2.180000  1.835000 3.135000 2.085000 ;
      RECT 2.180000  2.085000 2.510000 2.295000 ;
      RECT 2.210000  0.255000 3.595000 0.465000 ;
      RECT 2.210000  0.465000 2.540000 0.655000 ;
      RECT 2.710000  0.635000 3.135000 0.825000 ;
      RECT 2.965000  0.825000 3.135000 1.835000 ;
      RECT 3.305000  0.465000 3.595000 0.735000 ;
      RECT 3.305000  1.495000 3.595000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o32a_1
MACRO sky130_fd_sc_hd__o32a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495000 0.995000 1.715000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.995000 2.160000 1.615000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415000 0.995000 2.635000 1.615000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.695000 1.075000 4.055000 1.245000 ;
        RECT 3.725000 1.245000 4.055000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.910000 0.995000 3.155000 1.615000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.845000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.885000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 1.015000  0.995000 1.325000 1.785000 ;
      RECT 1.015000  1.785000 3.525000 1.955000 ;
      RECT 1.015000  2.125000 1.525000 2.635000 ;
      RECT 1.095000  0.085000 1.425000 0.825000 ;
      RECT 1.695000  0.255000 2.025000 0.655000 ;
      RECT 1.695000  0.655000 3.025000 0.825000 ;
      RECT 2.195000  0.085000 2.525000 0.485000 ;
      RECT 2.695000  0.255000 4.055000 0.425000 ;
      RECT 2.695000  0.425000 3.025000 0.655000 ;
      RECT 2.695000  1.955000 3.025000 2.465000 ;
      RECT 3.195000  0.595000 3.525000 0.825000 ;
      RECT 3.325000  0.825000 3.525000 1.785000 ;
      RECT 3.695000  0.425000 4.055000 0.905000 ;
      RECT 3.695000  1.495000 4.055000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__o32a_2
MACRO sky130_fd_sc_hd__o32a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 1.075000 0.780000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 1.075000 1.700000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.010000 1.075000 2.625000 1.275000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.870000 1.075000 4.230000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.790000 1.075000 5.260000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.305000 0.255000 6.635000 0.715000 ;
        RECT 6.305000 0.715000 8.135000 0.905000 ;
        RECT 6.305000 1.495000 8.135000 1.665000 ;
        RECT 6.305000 1.665000 6.635000 2.465000 ;
        RECT 7.145000 0.255000 7.475000 0.715000 ;
        RECT 7.145000 1.665000 7.475000 2.465000 ;
        RECT 7.645000 0.905000 8.135000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.635000 ;
      RECT 0.085000  0.635000 2.965000 0.885000 ;
      RECT 0.085000  1.445000 1.265000 1.665000 ;
      RECT 0.085000  1.665000 0.425000 2.465000 ;
      RECT 0.515000  0.085000 2.545000 0.465000 ;
      RECT 0.595000  1.835000 0.765000 2.635000 ;
      RECT 0.935000  1.665000 1.265000 2.295000 ;
      RECT 0.935000  2.295000 2.105000 2.465000 ;
      RECT 1.435000  1.445000 2.625000 1.690000 ;
      RECT 1.435000  1.690000 1.605000 2.045000 ;
      RECT 1.775000  1.860000 2.105000 2.295000 ;
      RECT 2.295000  1.690000 2.625000 2.295000 ;
      RECT 2.295000  2.295000 3.465000 2.465000 ;
      RECT 2.715000  0.255000 5.695000 0.465000 ;
      RECT 2.715000  0.465000 2.965000 0.635000 ;
      RECT 2.795000  1.105000 3.645000 1.275000 ;
      RECT 2.795000  1.275000 2.965000 2.045000 ;
      RECT 3.135000  1.445000 3.465000 2.295000 ;
      RECT 3.455000  0.635000 5.775000 0.805000 ;
      RECT 3.455000  0.805000 3.645000 1.105000 ;
      RECT 3.655000  1.445000 3.985000 1.785000 ;
      RECT 3.655000  1.785000 4.825000 1.955000 ;
      RECT 3.655000  1.955000 3.985000 2.465000 ;
      RECT 4.155000  2.125000 4.325000 2.635000 ;
      RECT 4.400000  0.805000 4.620000 1.445000 ;
      RECT 4.400000  1.445000 5.195000 1.615000 ;
      RECT 4.495000  1.955000 4.825000 2.285000 ;
      RECT 4.495000  2.285000 5.695000 2.465000 ;
      RECT 5.025000  1.615000 5.195000 2.115000 ;
      RECT 5.365000  1.445000 5.695000 2.285000 ;
      RECT 5.520000  0.805000 5.775000 1.075000 ;
      RECT 5.520000  1.075000 7.475000 1.245000 ;
      RECT 5.520000  1.245000 6.135000 1.265000 ;
      RECT 5.965000  0.085000 6.135000 0.885000 ;
      RECT 5.965000  1.835000 6.135000 2.635000 ;
      RECT 6.805000  0.085000 6.975000 0.545000 ;
      RECT 6.805000  1.835000 6.975000 2.635000 ;
      RECT 7.645000  0.085000 7.900000 0.545000 ;
      RECT 7.645000  1.835000 7.900000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
END sky130_fd_sc_hd__o32a_4
MACRO sky130_fd_sc_hd__o32ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.575000 0.995000 3.135000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.930000 0.995000 2.225000 2.465000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.410000 0.995000 1.700000 1.615000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.685000 0.345000 0.995000 ;
        RECT 0.090000 0.995000 0.360000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.870000 0.995000 1.240000 1.615000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.821250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.655000 0.845000 0.825000 ;
        RECT 0.530000 0.825000 0.700000 1.785000 ;
        RECT 0.530000 1.785000 1.545000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  0.255000 1.345000 0.485000 ;
      RECT 0.090000  1.495000 0.360000 2.635000 ;
      RECT 1.015000  0.485000 1.345000 0.655000 ;
      RECT 1.015000  0.655000 2.525000 0.825000 ;
      RECT 1.515000  0.085000 2.185000 0.485000 ;
      RECT 2.355000  0.375000 2.525000 0.655000 ;
      RECT 2.695000  0.085000 3.135000 0.825000 ;
      RECT 2.695000  1.495000 3.135000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o32ai_1
MACRO sky130_fd_sc_hd__o32ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.750000 1.075000 5.865000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.370000 1.075000 4.480000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 1.075000 3.065000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 1.075000 1.705000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.845000 1.325000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.655000 2.045000 0.905000 ;
        RECT 0.515000 1.495000 3.105000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.095000 ;
        RECT 1.875000 0.905000 2.045000 1.105000 ;
        RECT 1.875000 1.105000 2.170000 1.495000 ;
        RECT 2.775000 1.665000 3.105000 2.085000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.090000  0.255000 2.405000 0.485000 ;
      RECT 0.090000  0.485000 0.345000 0.905000 ;
      RECT 0.090000  1.495000 0.345000 2.295000 ;
      RECT 0.090000  2.295000 1.265000 2.465000 ;
      RECT 1.015000  1.835000 2.105000 2.005000 ;
      RECT 1.015000  2.005000 1.265000 2.295000 ;
      RECT 1.435000  2.175000 1.605000 2.635000 ;
      RECT 1.775000  2.005000 2.105000 2.455000 ;
      RECT 2.235000  0.485000 2.405000 0.715000 ;
      RECT 2.235000  0.715000 5.755000 0.905000 ;
      RECT 2.335000  1.835000 2.585000 2.255000 ;
      RECT 2.335000  2.255000 4.385000 2.445000 ;
      RECT 2.620000  0.085000 2.950000 0.545000 ;
      RECT 3.135000  0.255000 3.465000 0.715000 ;
      RECT 3.275000  1.495000 3.445000 2.255000 ;
      RECT 3.615000  1.495000 5.325000 1.665000 ;
      RECT 3.615000  1.665000 3.945000 2.085000 ;
      RECT 3.635000  0.085000 3.805000 0.545000 ;
      RECT 4.055000  0.255000 4.725000 0.715000 ;
      RECT 4.135000  1.835000 4.385000 2.255000 ;
      RECT 4.620000  1.835000 4.825000 2.635000 ;
      RECT 4.905000  0.085000 5.235000 0.545000 ;
      RECT 4.995000  1.665000 5.325000 2.460000 ;
      RECT 5.425000  0.255000 5.755000 0.715000 ;
      RECT 5.495000  1.495000 5.715000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__o32ai_2
MACRO sky130_fd_sc_hd__o32ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.290000 1.075000 10.035000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.090000 1.075000 7.260000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.770000 1.075000 5.380000 1.275000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.205000 1.075000 3.540000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 1.685000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.655000 3.380000 0.905000 ;
        RECT 0.515000 1.495000 5.580000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.085000 ;
        RECT 1.355000 1.665000 1.700000 2.085000 ;
        RECT 1.855000 0.905000 2.035000 1.495000 ;
        RECT 4.410000 1.665000 4.740000 2.085000 ;
        RECT 5.250000 1.665000 5.580000 2.085000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.090000  0.255000  3.800000 0.465000 ;
      RECT 0.090000  0.465000  0.345000 0.905000 ;
      RECT 0.090000  1.495000  0.345000 2.255000 ;
      RECT 0.090000  2.255000  2.040000 2.465000 ;
      RECT 1.015000  1.835000  1.185000 2.255000 ;
      RECT 1.870000  1.835000  3.800000 2.005000 ;
      RECT 1.870000  2.005000  2.040000 2.255000 ;
      RECT 2.210000  2.175000  2.540000 2.635000 ;
      RECT 2.710000  2.005000  2.880000 2.425000 ;
      RECT 3.050000  2.175000  3.380000 2.635000 ;
      RECT 3.550000  0.465000  3.800000 0.735000 ;
      RECT 3.550000  0.735000 10.035000 0.905000 ;
      RECT 3.550000  2.005000  3.800000 2.465000 ;
      RECT 3.970000  0.085000  4.140000 0.545000 ;
      RECT 3.990000  1.835000  4.240000 2.255000 ;
      RECT 3.990000  2.255000  7.680000 2.465000 ;
      RECT 4.310000  0.255000  4.640000 0.735000 ;
      RECT 4.810000  0.085000  5.140000 0.545000 ;
      RECT 4.910000  1.835000  5.080000 2.255000 ;
      RECT 5.310000  0.255000  5.980000 0.735000 ;
      RECT 5.750000  1.835000  5.920000 2.255000 ;
      RECT 6.090000  1.495000  9.460000 1.665000 ;
      RECT 6.090000  1.665000  6.420000 2.085000 ;
      RECT 6.170000  0.085000  6.340000 0.545000 ;
      RECT 6.510000  0.255000  6.840000 0.735000 ;
      RECT 6.590000  1.835000  6.760000 2.255000 ;
      RECT 6.930000  1.665000  7.260000 2.085000 ;
      RECT 7.010000  0.085000  7.180000 0.545000 ;
      RECT 7.350000  0.255000  8.040000 0.735000 ;
      RECT 7.430000  1.835000  7.680000 2.255000 ;
      RECT 7.870000  1.835000  8.120000 2.635000 ;
      RECT 8.290000  1.665000  8.620000 2.465000 ;
      RECT 8.370000  0.085000  8.540000 0.545000 ;
      RECT 8.710000  0.255000  9.040000 0.735000 ;
      RECT 8.790000  1.835000  8.960000 2.635000 ;
      RECT 9.130000  1.665000  9.460000 2.465000 ;
      RECT 9.210000  0.085000  9.470000 0.545000 ;
      RECT 9.630000  1.495000 10.035000 2.635000 ;
      RECT 9.645000  0.255000 10.035000 0.735000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
END sky130_fd_sc_hd__o32ai_4
MACRO sky130_fd_sc_hd__o41a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.075000 3.995000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 1.075000 3.275000 2.390000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 1.075000 2.735000 2.390000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.865000 1.075000 2.195000 2.390000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.275000 1.075000 1.695000 1.285000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.672000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.425000 0.885000 ;
        RECT 0.085000 0.885000 0.355000 1.455000 ;
        RECT 0.085000 1.455000 0.610000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.525000  1.075000 1.105000 1.285000 ;
      RECT 0.715000  0.085000 0.885000 0.545000 ;
      RECT 0.735000  0.715000 1.485000 0.905000 ;
      RECT 0.735000  0.905000 1.105000 1.075000 ;
      RECT 0.845000  1.285000 1.105000 1.455000 ;
      RECT 0.845000  1.455000 1.595000 1.745000 ;
      RECT 0.845000  1.915000 1.175000 2.635000 ;
      RECT 1.155000  0.270000 1.485000 0.715000 ;
      RECT 1.345000  1.745000 1.595000 2.465000 ;
      RECT 1.655000  0.415000 1.825000 0.735000 ;
      RECT 1.655000  0.735000 3.955000 0.905000 ;
      RECT 2.050000  0.085000 2.380000 0.545000 ;
      RECT 2.580000  0.255000 2.910000 0.735000 ;
      RECT 3.125000  0.085000 3.455000 0.545000 ;
      RECT 3.605000  1.515000 3.935000 2.635000 ;
      RECT 3.625000  0.255000 3.955000 0.735000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__o41a_1
MACRO sky130_fd_sc_hd__o41a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825000 1.075000 4.515000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.325000 1.075000 3.655000 2.335000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.825000 1.075000 3.155000 2.340000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 1.075000 2.655000 2.340000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775000 1.075000 2.155000 1.325000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.845000 0.880000 ;
        RECT 0.515000 0.880000 0.790000 1.495000 ;
        RECT 0.515000 1.495000 0.845000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.885000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 0.960000  1.075000 1.600000 1.325000 ;
      RECT 1.015000  0.085000 1.260000 0.885000 ;
      RECT 1.015000  1.495000 1.185000 1.835000 ;
      RECT 1.015000  1.835000 1.525000 2.635000 ;
      RECT 1.355000  1.325000 1.600000 1.495000 ;
      RECT 1.355000  1.495000 2.145000 1.665000 ;
      RECT 1.430000  0.255000 1.785000 0.850000 ;
      RECT 1.430000  0.850000 1.600000 1.075000 ;
      RECT 1.695000  1.665000 2.145000 2.465000 ;
      RECT 1.985000  0.255000 2.315000 0.715000 ;
      RECT 1.985000  0.715000 4.395000 0.905000 ;
      RECT 2.485000  0.085000 2.750000 0.545000 ;
      RECT 2.955000  0.255000 3.285000 0.715000 ;
      RECT 3.505000  0.085000 3.775000 0.545000 ;
      RECT 4.065000  0.255000 4.395000 0.715000 ;
      RECT 4.065000  1.495000 4.395000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__o41a_2
MACRO sky130_fd_sc_hd__o41a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.650000 1.075000 7.735000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.150000 1.075000 6.360000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.330000 1.075000 4.960000 1.275000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.410000 1.075000 4.040000 1.275000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.835000 1.075000 3.165000 1.275000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 1.685000 0.905000 ;
        RECT 0.085000 0.905000 0.345000 1.465000 ;
        RECT 0.085000 1.465000 1.685000 1.665000 ;
        RECT 0.515000 0.255000 0.845000 0.715000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 0.255000 1.685000 0.715000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.545000 ;
      RECT 0.085000  1.835000 0.345000 2.635000 ;
      RECT 0.515000  1.075000 2.665000 1.245000 ;
      RECT 0.515000  1.245000 2.545000 1.295000 ;
      RECT 1.015000  0.085000 1.185000 0.545000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.855000  0.085000 2.105000 0.885000 ;
      RECT 1.855000  1.465000 2.025000 2.635000 ;
      RECT 2.195000  1.295000 2.545000 1.445000 ;
      RECT 2.195000  1.445000 3.825000 1.615000 ;
      RECT 2.195000  1.615000 2.545000 2.465000 ;
      RECT 2.295000  0.255000 3.485000 0.465000 ;
      RECT 2.295000  0.635000 3.045000 0.905000 ;
      RECT 2.295000  0.905000 2.665000 1.075000 ;
      RECT 2.715000  1.835000 2.965000 2.635000 ;
      RECT 3.135000  1.835000 3.405000 2.295000 ;
      RECT 3.135000  2.295000 4.325000 2.465000 ;
      RECT 3.235000  0.465000 3.485000 0.735000 ;
      RECT 3.235000  0.735000 7.595000 0.905000 ;
      RECT 3.575000  1.615000 3.825000 2.125000 ;
      RECT 3.655000  0.085000 3.875000 0.545000 ;
      RECT 3.995000  1.445000 5.165000 1.615000 ;
      RECT 3.995000  1.615000 4.325000 2.295000 ;
      RECT 4.075000  0.255000 4.245000 0.735000 ;
      RECT 4.445000  0.085000 4.715000 0.545000 ;
      RECT 4.495000  1.785000 4.665000 2.295000 ;
      RECT 4.495000  2.295000 6.145000 2.465000 ;
      RECT 4.835000  1.615000 5.165000 2.115000 ;
      RECT 4.915000  0.255000 5.085000 0.735000 ;
      RECT 5.305000  0.085000 5.915000 0.545000 ;
      RECT 5.395000  1.445000 7.595000 1.615000 ;
      RECT 5.395000  1.615000 5.645000 2.115000 ;
      RECT 5.815000  1.785000 6.145000 2.295000 ;
      RECT 6.240000  0.255000 6.410000 0.735000 ;
      RECT 6.315000  1.615000 6.485000 2.455000 ;
      RECT 6.655000  1.785000 6.985000 2.635000 ;
      RECT 6.685000  0.085000 6.955000 0.545000 ;
      RECT 7.265000  0.255000 7.595000 0.735000 ;
      RECT 7.265000  1.615000 7.595000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__o41a_4
MACRO sky130_fd_sc_hd__o41ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.500000 1.075000 3.080000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 1.415000 2.330000 2.355000 ;
        RECT 2.000000 1.075000 2.330000 1.415000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 1.075000 1.830000 1.245000 ;
        RECT 1.500000 1.245000 1.820000 2.355000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.990000 1.075000 1.320000 1.245000 ;
        RECT 1.015000 1.245000 1.320000 2.355000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 0.440000 1.275000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.425000 0.735000 ;
        RECT 0.085000 0.735000 0.780000 0.905000 ;
        RECT 0.515000 1.485000 0.845000 2.465000 ;
        RECT 0.610000 0.905000 0.780000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  1.445000 0.345000 2.635000 ;
      RECT 0.790000  0.255000 1.120000 0.565000 ;
      RECT 0.950000  0.565000 1.120000 0.735000 ;
      RECT 0.950000  0.735000 2.960000 0.905000 ;
      RECT 1.290000  0.085000 1.540000 0.565000 ;
      RECT 1.710000  0.255000 2.040000 0.735000 ;
      RECT 2.210000  0.085000 2.460000 0.565000 ;
      RECT 2.630000  0.255000 2.960000 0.735000 ;
      RECT 2.630000  1.495000 2.960000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o41ai_1
MACRO sky130_fd_sc_hd__o41ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.720000 1.075000 5.895000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.780000 1.075000 4.540000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.595000 1.075000 3.580000 1.275000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 1.075000 2.325000 1.275000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 0.440000 1.275000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.635000 0.845000 0.885000 ;
        RECT 0.515000 1.505000 2.205000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 0.610000 0.885000 0.845000 1.445000 ;
        RECT 0.610000 1.445000 2.205000 1.505000 ;
        RECT 1.875000 1.665000 2.205000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.255000 1.265000 0.465000 ;
      RECT 0.085000  0.465000 0.345000 0.905000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 1.015000  0.465000 1.265000 0.735000 ;
      RECT 1.015000  0.735000 5.705000 0.905000 ;
      RECT 1.015000  1.835000 1.265000 2.635000 ;
      RECT 1.455000  0.085000 1.705000 0.545000 ;
      RECT 1.455000  1.835000 1.705000 2.295000 ;
      RECT 1.455000  2.295000 2.545000 2.465000 ;
      RECT 1.875000  0.255000 2.205000 0.735000 ;
      RECT 2.375000  0.085000 2.545000 0.545000 ;
      RECT 2.375000  1.445000 3.465000 1.615000 ;
      RECT 2.375000  1.615000 2.545000 2.295000 ;
      RECT 2.715000  0.255000 3.045000 0.735000 ;
      RECT 2.715000  1.835000 3.045000 2.295000 ;
      RECT 2.715000  2.295000 4.445000 2.465000 ;
      RECT 3.215000  0.085000 3.450000 0.545000 ;
      RECT 3.215000  1.615000 3.465000 2.125000 ;
      RECT 3.695000  0.255000 4.025000 0.735000 ;
      RECT 3.695000  1.445000 5.705000 1.615000 ;
      RECT 3.695000  1.615000 3.945000 2.125000 ;
      RECT 4.115000  1.835000 4.445000 2.295000 ;
      RECT 4.195000  0.085000 4.365000 0.545000 ;
      RECT 4.535000  0.255000 4.865000 0.735000 ;
      RECT 4.615000  1.615000 4.785000 2.465000 ;
      RECT 4.955000  1.785000 5.285000 2.635000 ;
      RECT 5.035000  0.085000 5.205000 0.545000 ;
      RECT 5.375000  0.255000 5.705000 0.735000 ;
      RECT 5.455000  1.615000 5.705000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__o41ai_2
MACRO sky130_fd_sc_hd__o41ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.155000 1.075000 10.035000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.170000 1.075000 7.940000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.310000 1.075000 5.980000 1.275000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.350000 1.075000 4.020000 1.275000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 1.700000 1.275000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.635000 2.160000 0.905000 ;
        RECT 0.515000 1.445000 3.885000 1.615000 ;
        RECT 0.515000 1.615000 0.845000 2.465000 ;
        RECT 1.355000 1.615000 1.685000 2.465000 ;
        RECT 1.870000 0.905000 2.160000 1.445000 ;
        RECT 2.715000 1.615000 3.045000 2.125000 ;
        RECT 3.555000 1.615000 3.885000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.085000  0.255000  2.625000 0.465000 ;
      RECT 0.085000  0.465000  0.345000 0.905000 ;
      RECT 0.085000  1.445000  0.345000 2.635000 ;
      RECT 1.015000  1.835000  1.185000 2.635000 ;
      RECT 1.855000  1.835000  2.105000 2.635000 ;
      RECT 2.295000  1.785000  2.545000 2.295000 ;
      RECT 2.295000  2.295000  4.225000 2.465000 ;
      RECT 2.350000  0.465000  2.625000 0.735000 ;
      RECT 2.350000  0.735000  9.865000 0.905000 ;
      RECT 2.795000  0.085000  2.965000 0.545000 ;
      RECT 3.135000  0.255000  3.465000 0.735000 ;
      RECT 3.215000  1.785000  3.385000 2.295000 ;
      RECT 3.635000  0.085000  3.805000 0.545000 ;
      RECT 3.975000  0.255000  4.305000 0.735000 ;
      RECT 4.055000  1.445000  5.985000 1.615000 ;
      RECT 4.055000  1.615000  4.225000 2.295000 ;
      RECT 4.395000  1.785000  4.645000 2.295000 ;
      RECT 4.395000  2.295000  7.685000 2.465000 ;
      RECT 4.475000  0.085000  4.645000 0.545000 ;
      RECT 4.815000  0.255000  5.145000 0.735000 ;
      RECT 4.815000  1.615000  5.145000 2.125000 ;
      RECT 5.315000  0.085000  5.485000 0.545000 ;
      RECT 5.315000  1.785000  5.485000 2.295000 ;
      RECT 5.655000  0.255000  5.985000 0.735000 ;
      RECT 5.655000  1.615000  5.985000 2.125000 ;
      RECT 6.175000  0.260000  6.505000 0.735000 ;
      RECT 6.175000  1.445000  9.865000 1.615000 ;
      RECT 6.175000  1.615000  6.505000 2.125000 ;
      RECT 6.675000  0.085000  6.845000 0.545000 ;
      RECT 6.675000  1.785000  6.845000 2.295000 ;
      RECT 7.015000  0.260000  7.345000 0.735000 ;
      RECT 7.015000  1.615000  7.345000 2.125000 ;
      RECT 7.515000  0.085000  7.685000 0.545000 ;
      RECT 7.515000  1.785000  7.685000 2.295000 ;
      RECT 7.855000  0.260000  8.185000 0.735000 ;
      RECT 7.855000  1.615000  8.185000 2.465000 ;
      RECT 8.355000  0.085000  8.525000 0.545000 ;
      RECT 8.355000  1.835000  8.525000 2.635000 ;
      RECT 8.695000  0.260000  9.025000 0.735000 ;
      RECT 8.695000  1.615000  9.025000 2.465000 ;
      RECT 9.195000  0.085000  9.365000 0.545000 ;
      RECT 9.195000  1.835000  9.365000 2.635000 ;
      RECT 9.535000  0.260000  9.865000 0.735000 ;
      RECT 9.535000  1.615000  9.865000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
END sky130_fd_sc_hd__o41ai_4
MACRO sky130_fd_sc_hd__o211a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.300000 1.075000 1.720000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.890000 1.075000 2.220000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.390000 1.075000 2.720000 1.275000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.245000 1.075000 3.595000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.425000 0.885000 ;
        RECT 0.085000 0.885000 0.260000 1.495000 ;
        RECT 0.085000 1.495000 0.425000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.430000  1.075000 1.125000 1.245000 ;
      RECT 0.595000  0.085000 0.845000 0.885000 ;
      RECT 0.595000  1.495000 0.765000 2.635000 ;
      RECT 0.955000  1.245000 1.125000 1.495000 ;
      RECT 0.955000  1.495000 3.390000 1.665000 ;
      RECT 1.035000  0.255000 1.365000 0.735000 ;
      RECT 1.035000  0.735000 2.260000 0.905000 ;
      RECT 1.035000  1.835000 1.285000 2.635000 ;
      RECT 1.535000  0.085000 1.760000 0.545000 ;
      RECT 1.930000  0.255000 2.260000 0.735000 ;
      RECT 1.930000  1.665000 2.260000 2.465000 ;
      RECT 2.560000  1.835000 2.890000 2.635000 ;
      RECT 2.890000  0.255000 3.390000 0.865000 ;
      RECT 2.890000  0.865000 3.060000 1.495000 ;
      RECT 3.060000  1.665000 3.390000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o211a_1
MACRO sky130_fd_sc_hd__o211a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 0.995000 2.325000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 0.995000 1.820000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.880000 0.995000 1.240000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.360000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.720000 0.255000 3.050000 0.615000 ;
        RECT 2.720000 0.615000 3.540000 0.785000 ;
        RECT 2.810000 1.905000 3.540000 2.075000 ;
        RECT 2.810000 2.075000 3.000000 2.465000 ;
        RECT 3.345000 0.785000 3.540000 1.905000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.090000  1.510000 2.665000 1.765000 ;
      RECT 0.090000  1.765000 0.355000 2.465000 ;
      RECT 0.095000  0.255000 0.430000 0.425000 ;
      RECT 0.095000  0.425000 0.710000 0.825000 ;
      RECT 0.525000  1.935000 0.855000 2.635000 ;
      RECT 0.530000  0.825000 0.710000 1.510000 ;
      RECT 0.880000  0.635000 2.150000 0.825000 ;
      RECT 1.025000  1.765000 1.695000 2.465000 ;
      RECT 1.390000  0.085000 1.725000 0.465000 ;
      RECT 2.200000  1.935000 2.630000 2.635000 ;
      RECT 2.315000  0.085000 2.550000 0.525000 ;
      RECT 2.495000  0.995000 3.175000 1.325000 ;
      RECT 2.495000  1.325000 2.665000 1.510000 ;
      RECT 3.170000  2.255000 3.500000 2.635000 ;
      RECT 3.220000  0.085000 3.550000 0.445000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o211a_2
MACRO sky130_fd_sc_hd__o211a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.490000 1.035000 4.845000 1.495000 ;
        RECT 4.490000 1.495000 6.290000 1.685000 ;
        RECT 5.890000 1.035000 6.290000 1.495000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.030000 1.035000 5.705000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.540000 0.995000 2.830000 1.445000 ;
        RECT 2.540000 1.445000 4.280000 1.685000 ;
        RECT 3.950000 1.035000 4.280000 1.445000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.055000 1.035000 3.740000 1.275000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.911000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.635000 1.605000 0.805000 ;
        RECT 0.085000 0.805000 0.365000 1.435000 ;
        RECT 0.085000 1.435000 2.030000 1.700000 ;
        RECT 0.595000 0.255000 0.765000 0.615000 ;
        RECT 0.595000 0.615000 1.605000 0.635000 ;
        RECT 0.980000 1.700000 1.160000 2.465000 ;
        RECT 1.435000 0.255000 1.605000 0.615000 ;
        RECT 1.840000 1.700000 2.030000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.480000  1.870000 0.810000 2.635000 ;
      RECT 0.535000  1.065000 2.370000 1.265000 ;
      RECT 0.935000  0.085000 1.265000 0.445000 ;
      RECT 1.340000  1.870000 1.670000 2.635000 ;
      RECT 1.775000  0.085000 2.140000 0.465000 ;
      RECT 2.200000  0.635000 3.520000 0.815000 ;
      RECT 2.200000  0.815000 2.370000 1.065000 ;
      RECT 2.200000  1.265000 2.370000 1.855000 ;
      RECT 2.200000  1.855000 5.485000 2.025000 ;
      RECT 2.200000  2.200000 2.530000 2.635000 ;
      RECT 2.330000  0.255000 4.500000 0.465000 ;
      RECT 2.700000  2.025000 3.060000 2.465000 ;
      RECT 3.285000  2.195000 3.615000 2.635000 ;
      RECT 3.785000  2.025000 4.120000 2.465000 ;
      RECT 4.170000  0.465000 4.500000 0.695000 ;
      RECT 4.170000  0.695000 6.345000 0.865000 ;
      RECT 4.290000  2.195000 4.555000 2.635000 ;
      RECT 4.670000  0.085000 4.985000 0.525000 ;
      RECT 5.155000  0.255000 5.485000 0.695000 ;
      RECT 5.155000  2.025000 5.485000 2.465000 ;
      RECT 5.655000  0.085000 5.845000 0.525000 ;
      RECT 6.015000  0.255000 6.345000 0.695000 ;
      RECT 6.015000  1.915000 6.345000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__o211a_4
MACRO sky130_fd_sc_hd__o211ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.395000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.995000 0.980000 1.325000 ;
        RECT 0.605000 1.325000 0.775000 2.250000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.300000 0.995000 1.795000 1.325000 ;
        RECT 1.470000 1.325000 1.795000 1.615000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.970000 1.075000 2.300000 1.615000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.418250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 1.595000 1.275000 1.815000 ;
        RECT 0.945000 1.815000 2.675000 2.045000 ;
        RECT 0.945000 2.045000 1.275000 2.445000 ;
        RECT 1.965000 0.255000 2.675000 0.845000 ;
        RECT 1.975000 2.045000 2.675000 2.465000 ;
        RECT 2.470000 0.845000 2.675000 1.815000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.095000  0.255000 0.425000 0.615000 ;
      RECT 0.095000  0.615000 1.455000 0.825000 ;
      RECT 0.095000  1.575000 0.425000 2.635000 ;
      RECT 0.595000  0.085000 0.925000 0.445000 ;
      RECT 1.125000  0.255000 1.455000 0.615000 ;
      RECT 1.445000  2.275000 1.775000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__o211ai_1
MACRO sky130_fd_sc_hd__o211ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.505000 1.075000 4.455000 1.245000 ;
        RECT 3.560000 1.245000 4.455000 1.295000 ;
        RECT 4.115000 0.765000 4.455000 1.075000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.365000 1.075000 3.335000 1.355000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.075000 1.905000 1.365000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.375000 1.970000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.022000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.670000 0.875000 1.540000 ;
        RECT 0.545000 1.540000 3.155000 1.710000 ;
        RECT 0.545000 1.710000 0.805000 2.465000 ;
        RECT 1.475000 1.710000 1.665000 2.465000 ;
        RECT 2.825000 1.710000 3.155000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.095000  0.255000 2.165000 0.445000 ;
      RECT 0.115000  2.175000 0.375000 2.635000 ;
      RECT 0.975000  1.915000 1.305000 2.635000 ;
      RECT 1.045000  0.445000 2.165000 0.465000 ;
      RECT 1.045000  0.465000 1.235000 0.890000 ;
      RECT 1.405000  0.635000 3.945000 0.845000 ;
      RECT 1.835000  1.915000 2.165000 2.635000 ;
      RECT 2.395000  0.085000 2.725000 0.445000 ;
      RECT 2.395000  2.100000 2.655000 2.295000 ;
      RECT 2.395000  2.295000 3.515000 2.465000 ;
      RECT 3.255000  0.085000 3.585000 0.445000 ;
      RECT 3.325000  1.525000 4.445000 1.695000 ;
      RECT 3.325000  1.695000 3.515000 2.295000 ;
      RECT 3.685000  1.865000 4.015000 2.635000 ;
      RECT 3.755000  0.515000 3.945000 0.635000 ;
      RECT 4.115000  0.085000 4.445000 0.445000 ;
      RECT 4.185000  1.695000 4.445000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__o211ai_2
MACRO sky130_fd_sc_hd__o211ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.400000 1.075000 1.410000 1.330000 ;
        RECT 0.965000 1.330000 1.410000 1.515000 ;
        RECT 0.965000 1.515000 3.630000 1.685000 ;
        RECT 3.350000 0.995000 3.630000 1.515000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.705000 1.075000 3.180000 1.345000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.800000 0.995000 4.975000 1.410000 ;
        RECT 4.260000 1.410000 4.975000 1.515000 ;
        RECT 4.260000 1.515000 7.000000 1.685000 ;
        RECT 6.830000 0.995000 7.000000 1.515000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.370000 1.075000 6.440000 1.345000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.001000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 1.855000 7.680000 2.025000 ;
        RECT 1.805000 2.025000 3.470000 2.105000 ;
        RECT 4.045000 2.025000 7.680000 2.105000 ;
        RECT 5.280000 0.270000 6.735000 0.450000 ;
        RECT 6.565000 0.450000 6.735000 0.655000 ;
        RECT 6.565000 0.655000 7.350000 0.825000 ;
        RECT 7.170000 0.825000 7.350000 1.340000 ;
        RECT 7.170000 1.340000 7.680000 1.855000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.090000  1.665000 0.385000 2.635000 ;
      RECT 0.155000  0.535000 0.355000 0.625000 ;
      RECT 0.155000  0.625000 1.240000 0.695000 ;
      RECT 0.155000  0.695000 3.835000 0.795000 ;
      RECT 0.155000  0.795000 3.130000 0.865000 ;
      RECT 0.155000  0.865000 1.795000 0.905000 ;
      RECT 0.525000  0.085000 0.855000 0.445000 ;
      RECT 0.555000  1.860000 0.775000 1.935000 ;
      RECT 0.555000  1.935000 1.635000 2.105000 ;
      RECT 0.555000  2.105000 0.775000 2.190000 ;
      RECT 0.955000  2.275000 1.285000 2.635000 ;
      RECT 1.025000  0.425000 1.240000 0.625000 ;
      RECT 1.455000  2.105000 1.635000 2.275000 ;
      RECT 1.455000  2.275000 3.435000 2.465000 ;
      RECT 1.465000  0.085000 1.635000 0.525000 ;
      RECT 1.775000  0.625000 3.835000 0.695000 ;
      RECT 2.245000  0.085000 2.575000 0.445000 ;
      RECT 3.105000  0.085000 3.435000 0.445000 ;
      RECT 3.605000  0.255000 4.920000 0.455000 ;
      RECT 3.605000  0.455000 3.835000 0.625000 ;
      RECT 3.615000  2.195000 3.885000 2.635000 ;
      RECT 4.005000  0.635000 6.170000 0.815000 ;
      RECT 4.435000  2.275000 4.765000 2.635000 ;
      RECT 5.280000  2.275000 5.610000 2.635000 ;
      RECT 6.120000  2.275000 6.455000 2.635000 ;
      RECT 6.980000  0.310000 7.680000 0.480000 ;
      RECT 7.355000  2.275000 7.685000 2.635000 ;
      RECT 7.510000  0.480000 7.680000 0.595000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  0.425000 1.240000 0.595000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.510000  0.425000 7.680000 0.595000 ;
    LAYER met1 ;
      RECT 1.010000 0.395000 1.300000 0.440000 ;
      RECT 1.010000 0.440000 7.740000 0.580000 ;
      RECT 1.010000 0.580000 1.300000 0.625000 ;
      RECT 7.450000 0.395000 7.740000 0.440000 ;
      RECT 7.450000 0.580000 7.740000 0.625000 ;
  END
END sky130_fd_sc_hd__o211ai_4
MACRO sky130_fd_sc_hd__o221a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.680000 1.075000 3.130000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005000 1.075000 2.490000 1.285000 ;
        RECT 2.005000 1.285000 2.380000 1.705000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.925000 1.075000 1.255000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 1.075000 1.815000 1.325000 ;
        RECT 1.495000 1.325000 1.815000 1.705000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.415000 1.285000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.370000 0.265000 4.055000 0.905000 ;
        RECT 3.390000 1.875000 4.055000 2.465000 ;
        RECT 3.805000 0.905000 4.055000 1.875000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.240000  1.455000 1.325000 1.625000 ;
      RECT 0.240000  1.625000 0.540000 2.465000 ;
      RECT 0.245000  0.255000 0.575000 0.645000 ;
      RECT 0.245000  0.645000 0.755000 0.825000 ;
      RECT 0.585000  0.825000 0.755000 1.455000 ;
      RECT 0.735000  1.795000 0.985000 2.635000 ;
      RECT 0.745000  0.305000 1.930000 0.475000 ;
      RECT 1.155000  1.625000 1.325000 1.875000 ;
      RECT 1.155000  1.875000 2.720000 2.045000 ;
      RECT 1.160000  0.645000 1.545000 0.735000 ;
      RECT 1.160000  0.735000 2.860000 0.905000 ;
      RECT 1.575000  2.045000 2.380000 2.465000 ;
      RECT 2.190000  0.085000 2.360000 0.555000 ;
      RECT 2.530000  0.270000 2.860000 0.735000 ;
      RECT 2.550000  1.455000 3.470000 1.625000 ;
      RECT 2.550000  1.625000 2.720000 1.875000 ;
      RECT 2.890000  1.795000 3.220000 2.635000 ;
      RECT 3.030000  0.085000 3.200000 0.905000 ;
      RECT 3.300000  1.075000 3.635000 1.285000 ;
      RECT 3.300000  1.285000 3.470000 1.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__o221a_1
MACRO sky130_fd_sc_hd__o221a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.635000 1.075000 3.075000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.980000 1.075000 2.465000 1.285000 ;
        RECT 1.980000 1.285000 2.285000 1.705000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.885000 1.075000 1.230000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.400000 1.075000 1.790000 1.275000 ;
        RECT 1.500000 1.275000 1.790000 1.705000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.345000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.295000 0.265000 3.625000 0.735000 ;
        RECT 3.295000 0.735000 4.055000 0.905000 ;
        RECT 3.295000 1.875000 4.055000 2.045000 ;
        RECT 3.295000 2.045000 3.545000 2.465000 ;
        RECT 3.745000 0.905000 4.055000 1.875000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.120000 -0.085000 0.290000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.170000  0.255000 0.500000 0.635000 ;
      RECT 0.170000  0.635000 0.715000 0.805000 ;
      RECT 0.250000  1.495000 1.330000 1.670000 ;
      RECT 0.250000  1.670000 0.580000 2.465000 ;
      RECT 0.545000  0.805000 0.715000 1.445000 ;
      RECT 0.545000  1.445000 1.330000 1.495000 ;
      RECT 0.670000  0.295000 1.855000 0.465000 ;
      RECT 0.750000  1.850000 0.990000 2.635000 ;
      RECT 1.085000  0.645000 1.470000 0.735000 ;
      RECT 1.085000  0.735000 2.785000 0.905000 ;
      RECT 1.160000  1.670000 1.330000 1.875000 ;
      RECT 1.160000  1.875000 2.625000 2.045000 ;
      RECT 1.550000  2.045000 2.305000 2.465000 ;
      RECT 2.115000  0.085000 2.285000 0.555000 ;
      RECT 2.455000  0.270000 2.785000 0.735000 ;
      RECT 2.455000  1.455000 3.415000 1.625000 ;
      RECT 2.455000  1.625000 2.625000 1.875000 ;
      RECT 2.795000  1.795000 3.125000 2.635000 ;
      RECT 2.955000  0.085000 3.125000 0.905000 ;
      RECT 3.245000  1.075000 3.575000 1.285000 ;
      RECT 3.245000  1.285000 3.415000 1.455000 ;
      RECT 3.715000  2.215000 4.055000 2.635000 ;
      RECT 3.795000  0.085000 3.965000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__o221a_2
MACRO sky130_fd_sc_hd__o221a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.075000 3.605000 1.445000 ;
        RECT 3.005000 1.445000 4.775000 1.615000 ;
        RECT 4.525000 1.075000 5.035000 1.275000 ;
        RECT 4.525000 1.275000 4.775000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775000 1.075000 4.355000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 1.075000 1.520000 1.445000 ;
        RECT 1.025000 1.445000 2.745000 1.615000 ;
        RECT 2.415000 1.075000 2.745000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.690000 1.075000 2.245000 1.275000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.440000 1.275000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235000 0.255000 5.565000 0.725000 ;
        RECT 5.235000 0.725000 6.405000 0.735000 ;
        RECT 5.235000 0.735000 6.920000 0.905000 ;
        RECT 5.315000 1.785000 5.900000 1.955000 ;
        RECT 5.315000 1.955000 5.525000 2.465000 ;
        RECT 5.730000 1.445000 6.920000 1.615000 ;
        RECT 5.730000 1.615000 5.900000 1.785000 ;
        RECT 6.075000 0.255000 6.405000 0.725000 ;
        RECT 6.115000 1.615000 6.365000 2.465000 ;
        RECT 6.575000 0.905000 6.920000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.085000  0.255000 2.955000 0.475000 ;
      RECT 0.085000  0.475000 0.345000 0.895000 ;
      RECT 0.145000  1.455000 0.395000 2.635000 ;
      RECT 0.515000  0.645000 0.845000 0.865000 ;
      RECT 0.565000  1.445000 0.845000 1.785000 ;
      RECT 0.565000  1.785000 5.145000 1.955000 ;
      RECT 0.565000  1.955000 0.815000 2.465000 ;
      RECT 0.610000  0.865000 0.845000 1.445000 ;
      RECT 0.985000  2.125000 1.235000 2.635000 ;
      RECT 1.015000  0.475000 1.185000 0.905000 ;
      RECT 1.355000  0.645000 2.535000 0.715000 ;
      RECT 1.355000  0.715000 3.885000 0.725000 ;
      RECT 1.355000  0.725000 4.725000 0.905000 ;
      RECT 1.405000  2.125000 1.655000 2.295000 ;
      RECT 1.405000  2.295000 2.495000 2.465000 ;
      RECT 1.825000  1.955000 2.075000 2.125000 ;
      RECT 2.245000  2.125000 2.495000 2.295000 ;
      RECT 2.665000  2.125000 3.425000 2.635000 ;
      RECT 3.145000  0.085000 3.385000 0.545000 ;
      RECT 3.555000  0.255000 3.885000 0.715000 ;
      RECT 3.595000  2.125000 3.845000 2.295000 ;
      RECT 3.595000  2.295000 4.685000 2.465000 ;
      RECT 4.015000  1.955000 4.265000 2.125000 ;
      RECT 4.055000  0.085000 4.225000 0.555000 ;
      RECT 4.395000  0.255000 4.725000 0.725000 ;
      RECT 4.435000  2.125000 4.685000 2.295000 ;
      RECT 4.855000  2.125000 5.105000 2.635000 ;
      RECT 4.895000  0.085000 5.065000 0.905000 ;
      RECT 4.975000  1.445000 5.375000 1.615000 ;
      RECT 4.975000  1.615000 5.145000 1.785000 ;
      RECT 5.205000  1.075000 6.405000 1.275000 ;
      RECT 5.205000  1.275000 5.375000 1.445000 ;
      RECT 5.695000  2.125000 5.945000 2.635000 ;
      RECT 5.735000  0.085000 5.905000 0.555000 ;
      RECT 6.535000  1.795000 6.785000 2.635000 ;
      RECT 6.575000  0.085000 6.830000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__o221a_4
MACRO sky130_fd_sc_hd__o221ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.675000 1.075000 3.135000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.165000 1.075000 2.505000 1.245000 ;
        RECT 2.295000 1.245000 2.505000 1.445000 ;
        RECT 2.295000 1.445000 2.675000 1.615000 ;
        RECT 2.465000 1.615000 2.675000 2.405000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.995000 1.355000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.995000 1.985000 1.325000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.465000 1.325000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.899000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.365000 0.345000 0.645000 ;
        RECT 0.085000 0.645000 0.840000 0.825000 ;
        RECT 0.085000 1.495000 2.125000 1.705000 ;
        RECT 0.085000 1.705000 0.365000 2.465000 ;
        RECT 0.635000 0.825000 0.840000 1.495000 ;
        RECT 1.735000 1.705000 2.125000 1.785000 ;
        RECT 1.735000 1.785000 2.245000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.515000  0.305000 1.775000 0.475000 ;
      RECT 0.550000  1.875000 1.340000 2.635000 ;
      RECT 1.010000  0.645000 2.220000 0.695000 ;
      RECT 1.010000  0.695000 3.135000 0.825000 ;
      RECT 1.945000  0.280000 2.220000 0.645000 ;
      RECT 2.105000  0.825000 3.135000 0.865000 ;
      RECT 2.455000  0.085000 2.625000 0.525000 ;
      RECT 2.795000  0.280000 3.135000 0.695000 ;
      RECT 2.875000  1.455000 3.135000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o221ai_1
MACRO sky130_fd_sc_hd__o221ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.430000 1.075000 3.760000 1.445000 ;
        RECT 3.430000 1.445000 4.815000 1.615000 ;
        RECT 4.645000 1.075000 5.435000 1.275000 ;
        RECT 4.645000 1.275000 4.815000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.980000 1.075000 4.475000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.020000 1.075000 2.035000 1.445000 ;
        RECT 1.020000 1.445000 3.260000 1.615000 ;
        RECT 2.930000 1.075000 3.260000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.205000 1.075000 2.760000 1.275000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.435000 1.275000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.985500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.520000 0.645000 0.850000 0.865000 ;
        RECT 0.560000 1.445000 0.850000 1.785000 ;
        RECT 0.560000 1.785000 4.350000 1.955000 ;
        RECT 0.560000 1.955000 0.810000 2.465000 ;
        RECT 0.605000 0.865000 0.850000 1.445000 ;
        RECT 2.340000 1.955000 2.590000 2.125000 ;
        RECT 4.100000 1.955000 4.350000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.100000  0.255000 1.270000 0.475000 ;
      RECT 0.100000  0.475000 0.350000 0.895000 ;
      RECT 0.140000  1.455000 0.390000 2.635000 ;
      RECT 0.980000  2.125000 1.750000 2.635000 ;
      RECT 1.020000  0.475000 1.270000 0.645000 ;
      RECT 1.020000  0.645000 3.050000 0.905000 ;
      RECT 1.460000  0.255000 3.550000 0.475000 ;
      RECT 1.920000  2.125000 2.170000 2.295000 ;
      RECT 1.920000  2.295000 3.010000 2.465000 ;
      RECT 2.760000  2.125000 3.010000 2.295000 ;
      RECT 3.180000  2.125000 3.510000 2.635000 ;
      RECT 3.220000  0.475000 3.550000 0.735000 ;
      RECT 3.220000  0.735000 5.230000 0.905000 ;
      RECT 3.680000  2.125000 3.930000 2.295000 ;
      RECT 3.680000  2.295000 4.770000 2.465000 ;
      RECT 3.720000  0.085000 3.890000 0.555000 ;
      RECT 4.060000  0.255000 4.390000 0.725000 ;
      RECT 4.060000  0.725000 5.230000 0.735000 ;
      RECT 4.520000  1.785000 4.770000 2.295000 ;
      RECT 4.560000  0.085000 4.730000 0.555000 ;
      RECT 4.900000  0.255000 5.230000 0.725000 ;
      RECT 4.985000  1.455000 5.190000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__o221ai_2
MACRO sky130_fd_sc_hd__o221ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.965000 1.075000 6.295000 1.445000 ;
        RECT 5.965000 1.445000 8.420000 1.615000 ;
        RECT 8.155000 1.075000 9.575000 1.275000 ;
        RECT 8.155000 1.275000 8.420000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.475000 1.075000 7.885000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.360000 1.075000 4.505000 1.275000 ;
        RECT 4.335000 1.275000 4.505000 1.495000 ;
        RECT 4.335000 1.495000 5.795000 1.665000 ;
        RECT 5.465000 1.075000 5.795000 1.495000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.675000 0.995000 5.285000 1.325000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.750000 1.275000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.971000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.645000 2.125000 0.865000 ;
        RECT 0.575000 1.445000 4.165000 1.615000 ;
        RECT 0.575000 1.615000 0.825000 2.465000 ;
        RECT 1.415000 1.615000 2.125000 1.955000 ;
        RECT 1.415000 1.955000 1.665000 2.465000 ;
        RECT 1.920000 0.865000 2.125000 1.445000 ;
        RECT 3.995000 1.615000 4.165000 1.835000 ;
        RECT 3.995000 1.835000 7.725000 1.955000 ;
        RECT 3.995000 1.955000 6.885000 2.005000 ;
        RECT 3.995000 2.005000 4.285000 2.125000 ;
        RECT 4.875000 2.005000 5.085000 2.125000 ;
        RECT 5.965000 1.785000 7.725000 1.835000 ;
        RECT 6.675000 2.005000 6.885000 2.125000 ;
        RECT 7.475000 1.955000 7.725000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.115000  0.255000 5.585000 0.475000 ;
      RECT 0.115000  0.475000 0.365000 0.895000 ;
      RECT 0.155000  1.485000 0.405000 2.635000 ;
      RECT 0.995000  1.825000 1.245000 2.635000 ;
      RECT 1.835000  2.125000 2.605000 2.635000 ;
      RECT 2.315000  0.645000 6.085000 0.735000 ;
      RECT 2.315000  0.735000 9.445000 0.820000 ;
      RECT 2.775000  1.785000 3.825000 1.955000 ;
      RECT 2.775000  1.955000 3.025000 2.465000 ;
      RECT 3.195000  2.125000 3.445000 2.635000 ;
      RECT 3.615000  1.955000 3.825000 2.295000 ;
      RECT 3.615000  2.295000 5.585000 2.465000 ;
      RECT 4.455000  2.175000 4.705000 2.295000 ;
      RECT 5.255000  2.175000 5.585000 2.295000 ;
      RECT 5.465000  0.820000 9.445000 0.905000 ;
      RECT 5.755000  0.255000 6.085000 0.645000 ;
      RECT 5.755000  2.175000 6.005000 2.635000 ;
      RECT 6.175000  2.175000 6.505000 2.295000 ;
      RECT 6.175000  2.295000 8.145000 2.465000 ;
      RECT 6.255000  0.085000 6.425000 0.555000 ;
      RECT 6.595000  0.255000 6.925000 0.725000 ;
      RECT 6.595000  0.725000 7.765000 0.735000 ;
      RECT 7.055000  2.125000 7.305000 2.295000 ;
      RECT 7.095000  0.085000 7.265000 0.555000 ;
      RECT 7.435000  0.255000 7.765000 0.725000 ;
      RECT 7.895000  1.785000 8.985000 1.955000 ;
      RECT 7.895000  1.955000 8.145000 2.295000 ;
      RECT 7.935000  0.085000 8.105000 0.555000 ;
      RECT 8.275000  0.255000 8.605000 0.725000 ;
      RECT 8.275000  0.725000 9.445000 0.735000 ;
      RECT 8.315000  2.125000 8.565000 2.635000 ;
      RECT 8.735000  1.445000 8.985000 1.785000 ;
      RECT 8.735000  1.955000 8.985000 2.465000 ;
      RECT 8.775000  0.085000 8.945000 0.555000 ;
      RECT 9.115000  0.255000 9.445000 0.725000 ;
      RECT 9.155000  1.445000 9.405000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
END sky130_fd_sc_hd__o221ai_4
MACRO sky130_fd_sc_hd__o311a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.995000 1.280000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.450000 0.995000 1.790000 1.325000 ;
        RECT 1.520000 1.325000 1.790000 2.070000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.980000 0.995000 2.270000 1.325000 ;
        RECT 1.980000 1.325000 2.215000 2.070000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.440000 0.995000 2.840000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.350000 0.995000 3.595000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.355000 1.070000 ;
        RECT 0.085000 1.070000 0.435000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.085000 0.310000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.525000  0.085000 1.195000 0.825000 ;
      RECT 0.605000  0.995000 0.775000 1.495000 ;
      RECT 0.605000  1.495000 1.350000 1.665000 ;
      RECT 0.605000  1.835000 1.010000 2.635000 ;
      RECT 1.180000  1.665000 1.350000 2.295000 ;
      RECT 1.180000  2.295000 2.715000 2.465000 ;
      RECT 1.365000  0.310000 1.660000 0.655000 ;
      RECT 1.365000  0.655000 2.760000 0.825000 ;
      RECT 1.840000  0.085000 2.215000 0.485000 ;
      RECT 2.385000  1.495000 3.595000 1.665000 ;
      RECT 2.385000  1.665000 2.715000 2.295000 ;
      RECT 2.430000  0.310000 2.760000 0.655000 ;
      RECT 2.900000  1.835000 3.135000 2.635000 ;
      RECT 3.010000  0.255000 3.595000 0.825000 ;
      RECT 3.010000  0.825000 3.180000 1.495000 ;
      RECT 3.305000  1.665000 3.595000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o311a_1
MACRO sky130_fd_sc_hd__o311a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 0.995000 1.750000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.920000 0.995000 2.250000 1.325000 ;
        RECT 1.980000 1.325000 2.250000 2.070000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.440000 0.995000 2.730000 1.325000 ;
        RECT 2.440000 1.325000 2.675000 2.070000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.900000 0.995000 3.300000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.810000 0.995000 4.055000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.905000 1.315000 ;
        RECT 0.550000 0.255000 0.825000 0.995000 ;
        RECT 0.550000 0.995000 0.905000 1.055000 ;
        RECT 0.550000 1.315000 0.905000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.085000 0.380000 0.885000 ;
      RECT 0.085000  1.485000 0.380000 2.635000 ;
      RECT 0.995000  0.085000 1.665000 0.825000 ;
      RECT 1.075000  0.995000 1.245000 1.495000 ;
      RECT 1.075000  1.495000 1.810000 1.665000 ;
      RECT 1.075000  1.835000 1.470000 2.635000 ;
      RECT 1.640000  1.665000 1.810000 2.295000 ;
      RECT 1.640000  2.295000 3.175000 2.465000 ;
      RECT 1.835000  0.310000 2.120000 0.655000 ;
      RECT 1.835000  0.655000 3.220000 0.825000 ;
      RECT 2.300000  0.085000 2.675000 0.485000 ;
      RECT 2.845000  1.495000 4.055000 1.665000 ;
      RECT 2.845000  1.665000 3.175000 2.295000 ;
      RECT 2.890000  0.310000 3.220000 0.655000 ;
      RECT 3.360000  1.835000 3.595000 2.635000 ;
      RECT 3.470000  0.255000 4.055000 0.825000 ;
      RECT 3.470000  0.825000 3.640000 1.495000 ;
      RECT 3.765000  1.665000 4.055000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__o311a_2
MACRO sky130_fd_sc_hd__o311a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.950000 1.055000 7.735000 1.315000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.020000 1.055000 6.770000 1.315000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.655000 1.055000 5.850000 1.315000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.250000 1.055000 4.475000 1.315000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.115000 1.055000 3.080000 1.315000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.765000 1.315000 ;
        RECT 0.595000 0.255000 0.765000 0.715000 ;
        RECT 0.595000 0.715000 1.605000 0.885000 ;
        RECT 0.595000 0.885000 0.765000 1.055000 ;
        RECT 0.595000 1.315000 0.765000 1.485000 ;
        RECT 0.595000 1.485000 1.605000 1.725000 ;
        RECT 0.595000 1.725000 0.765000 2.465000 ;
        RECT 1.435000 0.255000 1.605000 0.715000 ;
        RECT 1.435000 1.725000 1.605000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.085000  0.085000 0.425000 0.885000 ;
      RECT 0.085000  1.485000 0.425000 2.635000 ;
      RECT 0.935000  0.085000 1.265000 0.545000 ;
      RECT 0.935000  1.055000 1.945000 1.315000 ;
      RECT 0.935000  1.895000 1.265000 2.635000 ;
      RECT 1.775000  0.085000 2.025000 0.545000 ;
      RECT 1.775000  0.715000 3.045000 0.885000 ;
      RECT 1.775000  0.885000 1.945000 1.055000 ;
      RECT 1.775000  1.315000 1.945000 1.485000 ;
      RECT 1.775000  1.485000 5.005000 1.725000 ;
      RECT 1.775000  1.895000 2.445000 2.635000 ;
      RECT 2.195000  0.255000 4.305000 0.505000 ;
      RECT 2.195000  0.675000 3.045000 0.715000 ;
      RECT 2.615000  1.725000 2.785000 2.465000 ;
      RECT 2.955000  1.895000 3.285000 2.635000 ;
      RECT 3.215000  0.505000 3.385000 0.885000 ;
      RECT 3.455000  1.725000 3.625000 2.465000 ;
      RECT 3.555000  0.675000 7.735000 0.885000 ;
      RECT 3.855000  1.895000 4.045000 2.635000 ;
      RECT 4.335000  1.895000 4.665000 2.295000 ;
      RECT 4.335000  2.295000 6.445000 2.465000 ;
      RECT 4.485000  0.255000 4.755000 0.675000 ;
      RECT 4.835000  1.725000 5.005000 2.125000 ;
      RECT 4.925000  0.085000 5.605000 0.505000 ;
      RECT 5.255000  1.485000 5.525000 2.295000 ;
      RECT 5.695000  1.485000 7.735000 1.725000 ;
      RECT 5.695000  1.725000 5.945000 2.125000 ;
      RECT 5.775000  0.255000 5.945000 0.675000 ;
      RECT 6.115000  0.085000 6.445000 0.505000 ;
      RECT 6.115000  1.895000 6.445000 2.295000 ;
      RECT 6.615000  0.255000 6.785000 0.675000 ;
      RECT 6.615000  1.725000 6.785000 2.125000 ;
      RECT 6.955000  0.085000 7.285000 0.505000 ;
      RECT 6.955000  1.895000 7.285000 2.635000 ;
      RECT 7.455000  0.255000 7.735000 0.675000 ;
      RECT 7.455000  1.725000 7.735000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__o311a_4
MACRO sky130_fd_sc_hd__o311ai_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311ai_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.570000 0.995000 ;
        RECT 0.085000 0.995000 0.780000 1.625000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.995000 1.260000 2.465000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.430000 0.995000 1.780000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.260000 2.200000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.830000 0.765000 3.135000 1.325000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.604000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.430000 1.495000 3.135000 1.665000 ;
        RECT 1.430000 1.665000 1.980000 2.465000 ;
        RECT 2.445000 0.255000 3.135000 0.595000 ;
        RECT 2.445000 0.595000 2.660000 1.495000 ;
        RECT 2.650000 1.665000 3.135000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.085000 0.570000 0.595000 ;
      RECT 0.085000  1.795000 0.780000 2.635000 ;
      RECT 0.740000  0.255000 0.910000 0.655000 ;
      RECT 0.740000  0.655000 1.750000 0.825000 ;
      RECT 1.080000  0.085000 1.410000 0.485000 ;
      RECT 1.580000  0.255000 1.750000 0.655000 ;
      RECT 2.150000  1.835000 2.480000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o311ai_0
MACRO sky130_fd_sc_hd__o311ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.780000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.995000 1.260000 2.465000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.430000 0.995000 1.780000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.320000 2.200000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.830000 0.995000 3.135000 1.325000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.942000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.430000 1.495000 3.135000 1.665000 ;
        RECT 1.430000 1.665000 1.980000 2.465000 ;
        RECT 2.445000 0.255000 3.135000 0.825000 ;
        RECT 2.445000 0.825000 2.660000 1.495000 ;
        RECT 2.650000 1.665000 3.135000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.085000 0.570000 0.825000 ;
      RECT 0.085000  1.495000 0.780000 2.635000 ;
      RECT 0.740000  0.255000 0.910000 0.655000 ;
      RECT 0.740000  0.655000 1.750000 0.825000 ;
      RECT 1.080000  0.085000 1.410000 0.485000 ;
      RECT 1.580000  0.255000 1.750000 0.655000 ;
      RECT 2.150000  1.835000 2.480000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o311ai_1
MACRO sky130_fd_sc_hd__o311ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 1.105000 1.315000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.275000 1.055000 2.155000 1.315000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 1.055000 3.075000 1.315000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 1.055000 4.385000 1.315000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.085000 1.055000 5.895000 1.315000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.551000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415000 1.485000 5.895000 1.725000 ;
        RECT 2.415000 1.725000 2.665000 2.125000 ;
        RECT 3.335000 1.725000 3.505000 2.465000 ;
        RECT 4.515000 1.725000 4.825000 2.465000 ;
        RECT 4.555000 0.655000 5.895000 0.885000 ;
        RECT 4.555000 0.885000 4.915000 1.485000 ;
        RECT 5.495000 1.725000 5.895000 2.465000 ;
        RECT 5.515000 0.255000 5.895000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.255000 0.485000 0.655000 ;
      RECT 0.085000  0.655000 4.385000 0.885000 ;
      RECT 0.085000  1.485000 2.225000 1.725000 ;
      RECT 0.085000  1.725000 0.465000 2.465000 ;
      RECT 0.635000  1.895000 0.965000 2.635000 ;
      RECT 0.655000  0.085000 0.985000 0.485000 ;
      RECT 1.135000  1.725000 1.305000 2.465000 ;
      RECT 1.155000  0.255000 1.325000 0.655000 ;
      RECT 1.475000  1.895000 1.805000 2.295000 ;
      RECT 1.475000  2.295000 3.165000 2.465000 ;
      RECT 1.495000  0.085000 1.825000 0.485000 ;
      RECT 1.975000  1.725000 2.225000 2.125000 ;
      RECT 1.995000  0.255000 2.165000 0.655000 ;
      RECT 2.335000  0.085000 3.105000 0.485000 ;
      RECT 2.835000  1.895000 3.165000 2.295000 ;
      RECT 3.275000  0.255000 3.445000 0.655000 ;
      RECT 3.615000  0.255000 5.345000 0.485000 ;
      RECT 3.675000  1.895000 4.345000 2.635000 ;
      RECT 4.995000  1.895000 5.325000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__o311ai_2
MACRO sky130_fd_sc_hd__o311ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 1.775000 1.315000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 1.055000 3.615000 1.315000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 1.055000 5.885000 1.315000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.055000 1.055000 7.695000 1.315000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.865000 1.055000 9.090000 1.315000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.241000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.055000 1.485000 9.575000 1.725000 ;
        RECT 4.055000 1.725000 4.305000 2.115000 ;
        RECT 4.975000 1.725000 5.145000 2.115000 ;
        RECT 5.815000 1.725000 6.005000 2.465000 ;
        RECT 6.675000 1.725000 6.845000 2.465000 ;
        RECT 7.515000 1.725000 7.685000 2.465000 ;
        RECT 7.895000 0.655000 9.575000 0.885000 ;
        RECT 8.355000 1.725000 8.525000 2.465000 ;
        RECT 9.195000 1.725000 9.575000 2.465000 ;
        RECT 9.260000 0.885000 9.575000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.125000 -0.085000 0.295000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.085000  0.085000 0.505000 0.885000 ;
      RECT 0.085000  1.485000 3.865000 1.725000 ;
      RECT 0.085000  1.725000 0.405000 2.465000 ;
      RECT 0.595000  1.895000 0.925000 2.635000 ;
      RECT 0.675000  0.255000 0.845000 0.655000 ;
      RECT 0.675000  0.655000 7.385000 0.885000 ;
      RECT 1.015000  0.085000 1.345000 0.485000 ;
      RECT 1.095000  1.725000 1.265000 2.465000 ;
      RECT 1.435000  1.895000 1.765000 2.635000 ;
      RECT 1.515000  0.255000 1.685000 0.655000 ;
      RECT 1.855000  0.085000 2.185000 0.485000 ;
      RECT 1.935000  1.725000 2.105000 2.465000 ;
      RECT 2.275000  1.895000 2.605000 2.295000 ;
      RECT 2.275000  2.295000 5.645000 2.465000 ;
      RECT 2.355000  0.255000 2.525000 0.655000 ;
      RECT 2.695000  0.085000 3.025000 0.485000 ;
      RECT 2.775000  1.725000 2.945000 2.115000 ;
      RECT 3.115000  1.895000 3.445000 2.295000 ;
      RECT 3.195000  0.255000 3.365000 0.655000 ;
      RECT 3.535000  0.085000 3.885000 0.485000 ;
      RECT 3.615000  1.725000 3.865000 2.115000 ;
      RECT 4.055000  0.255000 4.225000 0.655000 ;
      RECT 4.395000  0.085000 4.725000 0.485000 ;
      RECT 4.475000  1.895000 4.805000 2.295000 ;
      RECT 4.895000  0.255000 5.065000 0.655000 ;
      RECT 5.235000  0.085000 5.585000 0.485000 ;
      RECT 5.315000  1.895000 5.645000 2.295000 ;
      RECT 5.755000  0.255000 9.575000 0.485000 ;
      RECT 6.175000  1.895000 6.505000 2.635000 ;
      RECT 7.015000  1.895000 7.345000 2.635000 ;
      RECT 7.555000  0.485000 7.725000 0.885000 ;
      RECT 7.855000  1.895000 8.185000 2.635000 ;
      RECT 8.695000  1.895000 9.025000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
END sky130_fd_sc_hd__o311ai_4
MACRO sky130_fd_sc_hd__o2111a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.705000 1.075000 4.035000 1.660000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.050000 1.075000 3.535000 1.325000 ;
        RECT 3.350000 1.325000 3.535000 2.415000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 0.390000 2.690000 0.995000 ;
        RECT 2.445000 0.995000 2.705000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925000 0.390000 2.195000 1.325000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.265000 1.075000 1.745000 1.325000 ;
        RECT 1.535000 0.390000 1.745000 1.075000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.255000 0.355000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.525000  0.995000 0.865000 1.325000 ;
      RECT 0.525000  1.835000 1.335000 2.635000 ;
      RECT 0.535000  0.085000 0.845000 0.565000 ;
      RECT 0.695000  0.735000 1.365000 0.905000 ;
      RECT 0.695000  0.905000 0.865000 0.995000 ;
      RECT 0.695000  1.325000 0.865000 1.495000 ;
      RECT 0.695000  1.495000 3.180000 1.665000 ;
      RECT 1.025000  0.255000 1.365000 0.735000 ;
      RECT 1.505000  1.665000 1.835000 2.465000 ;
      RECT 2.020000  1.835000 2.760000 2.635000 ;
      RECT 2.870000  0.255000 3.160000 0.705000 ;
      RECT 2.870000  0.705000 4.055000 0.875000 ;
      RECT 2.930000  1.665000 3.180000 2.465000 ;
      RECT 3.330000  0.085000 3.620000 0.535000 ;
      RECT 3.730000  1.835000 4.055000 2.635000 ;
      RECT 3.790000  0.255000 4.055000 0.705000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__o2111a_1
MACRO sky130_fd_sc_hd__o2111a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.830000 1.005000 4.515000 1.315000 ;
        RECT 4.310000 1.315000 4.515000 2.355000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.300000 0.995000 3.660000 1.325000 ;
        RECT 3.370000 1.325000 3.660000 2.370000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.680000 1.075000 3.100000 1.615000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005000 0.255000 2.390000 1.615000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.075000 1.835000 1.615000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.855000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.135000  0.085000 0.345000 0.885000 ;
      RECT 0.135000  1.495000 0.345000 2.635000 ;
      RECT 1.030000  0.715000 1.805000 0.885000 ;
      RECT 1.030000  0.885000 1.305000 1.785000 ;
      RECT 1.030000  1.785000 3.195000 2.025000 ;
      RECT 1.035000  0.085000 1.285000 0.545000 ;
      RECT 1.035000  2.195000 1.655000 2.635000 ;
      RECT 1.475000  0.255000 1.805000 0.715000 ;
      RECT 1.860000  2.025000 2.140000 2.465000 ;
      RECT 2.325000  2.255000 2.655000 2.635000 ;
      RECT 2.865000  0.255000 3.195000 0.625000 ;
      RECT 2.865000  0.625000 4.215000 0.825000 ;
      RECT 2.865000  2.025000 3.195000 2.465000 ;
      RECT 3.385000  0.085000 3.715000 0.455000 ;
      RECT 3.885000  0.255000 4.215000 0.625000 ;
      RECT 3.885000  1.495000 4.140000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__o2111a_2
MACRO sky130_fd_sc_hd__o2111a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.890000 1.075000 4.485000 1.245000 ;
        RECT 4.130000 1.245000 4.485000 1.320000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.135000 1.075000 3.600000 1.245000 ;
        RECT 3.145000 1.245000 3.600000 1.320000 ;
        RECT 3.305000 1.320000 3.600000 1.490000 ;
        RECT 3.305000 1.490000 4.825000 1.660000 ;
        RECT 4.655000 1.075000 4.985000 1.320000 ;
        RECT 4.655000 1.320000 4.825000 1.490000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775000 1.075000 2.215000 1.320000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.150000 0.995000 1.395000 1.490000 ;
        RECT 1.150000 1.490000 2.660000 1.660000 ;
        RECT 2.445000 1.080000 2.820000 1.320000 ;
        RECT 2.445000 1.320000 2.660000 1.490000 ;
        RECT 2.490000 1.075000 2.820000 1.080000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.995000 0.340000 1.655000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.962500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.650000 0.255000 5.875000 0.695000 ;
        RECT 5.650000 0.695000 7.275000 0.865000 ;
        RECT 5.755000 1.495000 7.275000 1.665000 ;
        RECT 5.755000 1.665000 5.925000 2.465000 ;
        RECT 6.545000 0.255000 6.745000 0.695000 ;
        RECT 6.585000 1.665000 6.775000 2.465000 ;
        RECT 7.005000 0.865000 7.275000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.090000  1.835000 5.550000 2.000000 ;
      RECT 0.090000  2.000000 5.065000 2.005000 ;
      RECT 0.090000  2.005000 0.345000 2.465000 ;
      RECT 0.100000  0.255000 2.940000 0.485000 ;
      RECT 0.100000  0.485000 0.345000 0.825000 ;
      RECT 0.515000  0.655000 0.860000 1.830000 ;
      RECT 0.515000  1.830000 5.550000 1.835000 ;
      RECT 0.515000  2.175000 0.845000 2.635000 ;
      RECT 1.015000  2.005000 1.230000 2.465000 ;
      RECT 1.400000  2.175000 1.625000 2.635000 ;
      RECT 1.720000  0.655000 4.795000 0.885000 ;
      RECT 1.795000  2.005000 2.025000 2.465000 ;
      RECT 2.195000  2.175000 2.525000 2.635000 ;
      RECT 2.695000  2.005000 3.285000 2.465000 ;
      RECT 3.110000  0.085000 3.440000 0.485000 ;
      RECT 3.610000  0.255000 3.825000 0.655000 ;
      RECT 3.805000  2.180000 4.135000 2.635000 ;
      RECT 3.995000  0.085000 4.365000 0.485000 ;
      RECT 4.535000  0.255000 4.795000 0.655000 ;
      RECT 4.775000  2.005000 5.065000 2.465000 ;
      RECT 5.035000  0.085000 5.300000 0.545000 ;
      RECT 5.245000  2.170000 5.585000 2.635000 ;
      RECT 5.380000  1.075000 6.760000 1.320000 ;
      RECT 5.380000  1.320000 5.550000 1.830000 ;
      RECT 6.075000  0.085000 6.375000 0.525000 ;
      RECT 6.095000  1.835000 6.415000 2.635000 ;
      RECT 6.915000  0.085000 7.275000 0.525000 ;
      RECT 6.945000  1.835000 7.270000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__o2111a_4
MACRO sky130_fd_sc_hd__o2111ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 1.005000 3.115000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.995000 2.615000 1.615000 ;
        RECT 2.270000 1.615000 2.615000 2.370000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.995000 1.815000 1.615000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 0.255000 1.355000 1.615000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.485000 1.075000 0.815000 1.615000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  0.857250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.690000 0.885000 ;
        RECT 0.085000 0.885000 0.315000 1.785000 ;
        RECT 0.085000 1.785000 2.095000 2.025000 ;
        RECT 0.790000 2.025000 1.025000 2.465000 ;
        RECT 1.750000 2.025000 2.095000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.290000  2.195000 0.620000 2.635000 ;
      RECT 1.210000  2.255000 1.540000 2.635000 ;
      RECT 1.750000  0.255000 2.095000 0.625000 ;
      RECT 1.750000  0.625000 3.115000 0.825000 ;
      RECT 2.285000  0.085000 2.615000 0.455000 ;
      RECT 2.785000  0.255000 3.115000 0.625000 ;
      RECT 2.785000  1.795000 3.115000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o2111ai_1
MACRO sky130_fd_sc_hd__o2111ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.635000 1.075000 5.435000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 1.075000 4.455000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.200000 1.075000 3.185000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.075000 1.790000 1.325000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.355000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.302000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.615000 0.935000 0.905000 ;
        RECT 0.605000 0.905000 0.865000 1.495000 ;
        RECT 0.605000 1.495000 4.005000 1.665000 ;
        RECT 0.605000 1.665000 0.865000 2.465000 ;
        RECT 1.535000 1.665000 1.725000 2.465000 ;
        RECT 2.395000 1.665000 2.575000 2.465000 ;
        RECT 3.815000 1.665000 4.005000 2.105000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.175000  0.260000 1.300000 0.445000 ;
      RECT 0.175000  0.445000 0.435000 0.865000 ;
      RECT 0.175000  1.525000 0.425000 2.635000 ;
      RECT 1.035000  1.835000 1.365000 2.635000 ;
      RECT 1.115000  0.445000 1.300000 0.735000 ;
      RECT 1.115000  0.735000 2.275000 0.905000 ;
      RECT 1.470000  0.255000 3.210000 0.445000 ;
      RECT 1.470000  0.445000 1.775000 0.530000 ;
      RECT 1.470000  0.530000 1.760000 0.565000 ;
      RECT 1.895000  1.840000 2.225000 2.635000 ;
      RECT 1.925000  0.620000 2.275000 0.735000 ;
      RECT 2.450000  0.655000 5.435000 0.840000 ;
      RECT 2.755000  1.835000 3.085000 2.635000 ;
      RECT 2.880000  0.445000 3.210000 0.485000 ;
      RECT 3.310000  1.835000 3.570000 2.275000 ;
      RECT 3.310000  2.275000 4.500000 2.465000 ;
      RECT 3.380000  0.365000 3.570000 0.655000 ;
      RECT 3.740000  0.085000 4.070000 0.485000 ;
      RECT 4.240000  0.365000 4.430000 0.650000 ;
      RECT 4.240000  0.650000 5.435000 0.655000 ;
      RECT 4.240000  1.515000 5.360000 1.685000 ;
      RECT 4.240000  1.685000 4.500000 2.275000 ;
      RECT 4.600000  0.085000 4.930000 0.480000 ;
      RECT 4.670000  1.855000 4.930000 2.635000 ;
      RECT 5.100000  0.365000 5.435000 0.650000 ;
      RECT 5.100000  1.685000 5.360000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__o2111ai_2
MACRO sky130_fd_sc_hd__o2111ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.820000 1.075000 9.575000 1.340000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.110000 1.075000 7.325000 1.345000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 1.075000 5.455000 1.345000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.940000 1.075000 3.550000 1.345000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.075000 1.755000 1.345000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  2.984350 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.645000 1.685000 0.815000 ;
        RECT 0.085000 0.815000 0.375000 1.515000 ;
        RECT 0.085000 1.515000 7.390000 1.685000 ;
        RECT 0.085000 1.685000 0.360000 2.465000 ;
        RECT 1.015000 1.685000 1.195000 2.465000 ;
        RECT 1.845000 1.685000 2.035000 2.465000 ;
        RECT 2.685000 1.685000 2.875000 2.465000 ;
        RECT 3.525000 1.685000 3.715000 2.465000 ;
        RECT 4.570000 1.685000 4.760000 2.465000 ;
        RECT 5.410000 1.685000 5.600000 2.465000 ;
        RECT 6.285000 1.685000 6.480000 2.100000 ;
        RECT 7.045000 1.685000 7.390000 1.720000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.095000  0.285000 2.025000 0.475000 ;
      RECT 0.530000  1.855000 0.845000 2.635000 ;
      RECT 1.390000  1.855000 1.675000 2.635000 ;
      RECT 1.855000  0.475000 2.025000 0.615000 ;
      RECT 1.855000  0.615000 3.785000 0.825000 ;
      RECT 2.195000  0.255000 5.565000 0.445000 ;
      RECT 2.205000  1.855000 2.515000 2.635000 ;
      RECT 3.045000  1.855000 3.355000 2.635000 ;
      RECT 3.975000  0.655000 9.440000 0.905000 ;
      RECT 4.075000  1.855000 4.400000 2.635000 ;
      RECT 4.930000  1.855000 5.220000 2.635000 ;
      RECT 5.785000  1.855000 6.115000 2.270000 ;
      RECT 5.785000  2.270000 7.005000 2.465000 ;
      RECT 6.100000  0.085000 6.430000 0.485000 ;
      RECT 6.705000  1.890000 8.235000 2.060000 ;
      RECT 6.705000  2.060000 7.005000 2.270000 ;
      RECT 6.960000  0.085000 7.290000 0.485000 ;
      RECT 7.555000  2.230000 7.885000 2.635000 ;
      RECT 7.825000  0.085000 8.155000 0.485000 ;
      RECT 8.045000  1.515000 9.080000 1.685000 ;
      RECT 8.045000  1.685000 8.235000 1.890000 ;
      RECT 8.055000  2.060000 8.235000 2.465000 ;
      RECT 8.410000  1.855000 8.720000 2.635000 ;
      RECT 8.665000  0.085000 8.995000 0.485000 ;
      RECT 8.890000  1.685000 9.080000 2.465000 ;
      RECT 9.265000  1.535000 9.575000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
END sky130_fd_sc_hd__o2111ai_4
MACRO sky130_fd_sc_hd__or2_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.995000 1.335000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.995000 0.500000 1.615000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.326800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.525000 2.180000 0.825000 ;
        RECT 1.645000 2.135000 2.180000 2.465000 ;
        RECT 1.865000 0.825000 2.180000 2.135000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.250000  0.085000 0.490000 0.825000 ;
      RECT 0.270000  1.785000 1.695000 1.955000 ;
      RECT 0.270000  1.955000 0.660000 2.130000 ;
      RECT 0.670000  0.425000 0.950000 0.825000 ;
      RECT 0.670000  0.825000 0.840000 1.785000 ;
      RECT 1.145000  2.125000 1.475000 2.635000 ;
      RECT 1.180000  0.085000 1.395000 0.825000 ;
      RECT 1.525000  0.995000 1.695000 1.785000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__or2_0
MACRO sky130_fd_sc_hd__or2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.765000 1.275000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.765000 0.500000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.509000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.255000 2.180000 0.825000 ;
        RECT 1.645000 1.845000 2.180000 2.465000 ;
        RECT 1.865000 0.825000 2.180000 1.845000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.250000  0.085000 0.490000 0.595000 ;
      RECT 0.270000  1.495000 1.695000 1.665000 ;
      RECT 0.270000  1.665000 0.660000 1.840000 ;
      RECT 0.670000  0.265000 0.950000 0.595000 ;
      RECT 0.670000  0.595000 0.840000 1.495000 ;
      RECT 1.145000  1.835000 1.475000 2.635000 ;
      RECT 1.180000  0.085000 1.395000 0.595000 ;
      RECT 1.525000  0.995000 1.695000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__or2_1
MACRO sky130_fd_sc_hd__or2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 0.765000 1.275000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.765000 0.345000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.440000 1.835000 2.215000 2.005000 ;
        RECT 1.440000 2.005000 1.770000 2.465000 ;
        RECT 1.520000 0.385000 1.690000 0.655000 ;
        RECT 1.520000 0.655000 2.215000 0.825000 ;
        RECT 1.785000 0.825000 2.215000 1.835000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.105000  0.085000 0.345000 0.595000 ;
      RECT 0.155000  1.495000 1.615000 1.665000 ;
      RECT 0.155000  1.665000 0.515000 1.840000 ;
      RECT 0.515000  0.255000 0.805000 0.595000 ;
      RECT 0.515000  0.595000 0.695000 1.495000 ;
      RECT 1.035000  0.085000 1.350000 0.595000 ;
      RECT 1.100000  1.835000 1.270000 2.635000 ;
      RECT 1.445000  0.995000 1.615000 1.495000 ;
      RECT 1.860000  0.085000 2.190000 0.485000 ;
      RECT 1.940000  2.175000 2.110000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__or2_2
MACRO sky130_fd_sc_hd__or2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 0.995000 1.240000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.765000 0.345000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.440000 0.265000 1.770000 0.735000 ;
        RECT 1.440000 0.735000 3.135000 0.905000 ;
        RECT 1.440000 1.835000 2.610000 2.005000 ;
        RECT 1.440000 2.005000 1.770000 2.465000 ;
        RECT 2.280000 0.265000 2.610000 0.735000 ;
        RECT 2.280000 1.495000 3.135000 1.665000 ;
        RECT 2.280000 1.665000 2.610000 1.835000 ;
        RECT 2.280000 2.005000 2.610000 2.465000 ;
        RECT 2.790000 0.905000 3.135000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.105000  0.085000 0.345000 0.595000 ;
      RECT 0.155000  1.495000 1.615000 1.665000 ;
      RECT 0.155000  1.665000 0.515000 2.465000 ;
      RECT 0.515000  0.290000 0.845000 0.825000 ;
      RECT 0.515000  0.825000 0.695000 1.495000 ;
      RECT 1.060000  0.085000 1.230000 0.825000 ;
      RECT 1.060000  1.835000 1.230000 2.635000 ;
      RECT 1.410000  1.075000 2.620000 1.245000 ;
      RECT 1.410000  1.245000 1.615000 1.495000 ;
      RECT 1.940000  0.085000 2.110000 0.565000 ;
      RECT 1.940000  2.175000 2.110000 2.635000 ;
      RECT 2.780000  0.085000 2.950000 0.565000 ;
      RECT 2.780000  1.835000 2.950000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__or2_4
MACRO sky130_fd_sc_hd__or2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 2.085000 1.735000 2.415000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.425000 1.325000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 0.415000 2.675000 0.760000 ;
        RECT 2.405000 1.495000 2.675000 2.465000 ;
        RECT 2.505000 0.760000 2.675000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.110000  0.265000 0.420000 0.735000 ;
      RECT 0.110000  0.735000 0.845000 0.905000 ;
      RECT 0.590000  0.085000 1.325000 0.565000 ;
      RECT 0.595000  0.905000 0.845000 0.995000 ;
      RECT 0.595000  0.995000 1.335000 1.325000 ;
      RECT 0.595000  1.325000 0.765000 1.885000 ;
      RECT 0.990000  1.495000 2.235000 1.665000 ;
      RECT 0.990000  1.665000 1.410000 1.915000 ;
      RECT 1.495000  0.305000 1.665000 0.655000 ;
      RECT 1.495000  0.655000 2.235000 0.825000 ;
      RECT 1.835000  0.085000 2.215000 0.485000 ;
      RECT 1.915000  1.835000 2.195000 2.635000 ;
      RECT 2.065000  0.825000 2.235000 0.995000 ;
      RECT 2.065000  0.995000 2.295000 1.325000 ;
      RECT 2.065000  1.325000 2.235000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__or2b_1
MACRO sky130_fd_sc_hd__or2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 2.085000 1.730000 2.415000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.325000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.400000 0.415000 2.630000 0.760000 ;
        RECT 2.400000 1.495000 2.630000 2.465000 ;
        RECT 2.460000 0.760000 2.630000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 0.105000  0.265000 0.420000 0.735000 ;
      RECT 0.105000  0.735000 0.840000 0.905000 ;
      RECT 0.590000  0.085000 1.320000 0.565000 ;
      RECT 0.595000  0.905000 0.840000 0.995000 ;
      RECT 0.595000  0.995000 1.330000 1.325000 ;
      RECT 0.595000  1.325000 0.765000 1.885000 ;
      RECT 0.985000  1.495000 2.230000 1.665000 ;
      RECT 0.985000  1.665000 1.405000 1.915000 ;
      RECT 1.490000  0.305000 1.660000 0.655000 ;
      RECT 1.490000  0.655000 2.230000 0.825000 ;
      RECT 1.830000  0.085000 2.210000 0.485000 ;
      RECT 1.910000  1.835000 2.190000 2.635000 ;
      RECT 2.060000  0.825000 2.230000 0.995000 ;
      RECT 2.060000  0.995000 2.290000 1.325000 ;
      RECT 2.060000  1.325000 2.230000 1.495000 ;
      RECT 2.800000  0.085000 3.055000 0.925000 ;
      RECT 2.800000  1.460000 3.055000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__or2b_2
MACRO sky130_fd_sc_hd__or2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.630000 1.075000 2.320000 1.275000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.425000 1.955000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 0.290000 2.655000 0.735000 ;
        RECT 2.325000 0.735000 4.055000 0.905000 ;
        RECT 2.365000 1.785000 3.455000 1.955000 ;
        RECT 2.365000 1.955000 2.615000 2.465000 ;
        RECT 2.830000 1.445000 4.055000 1.615000 ;
        RECT 2.830000 1.615000 3.455000 1.785000 ;
        RECT 3.165000 0.290000 3.495000 0.735000 ;
        RECT 3.205000 1.955000 3.455000 2.465000 ;
        RECT 3.670000 0.905000 4.055000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  2.125000 0.345000 2.635000 ;
      RECT 0.110000  0.265000 0.420000 0.735000 ;
      RECT 0.110000  0.735000 0.845000 0.905000 ;
      RECT 0.590000  0.085000 1.245000 0.565000 ;
      RECT 0.595000  0.905000 0.845000 0.995000 ;
      RECT 0.595000  0.995000 1.120000 1.325000 ;
      RECT 0.595000  1.325000 0.765000 2.465000 ;
      RECT 0.990000  1.495000 2.660000 1.615000 ;
      RECT 0.990000  1.615000 1.460000 2.465000 ;
      RECT 1.290000  0.735000 1.745000 0.905000 ;
      RECT 1.290000  0.905000 1.460000 1.445000 ;
      RECT 1.290000  1.445000 2.660000 1.495000 ;
      RECT 1.415000  0.305000 1.745000 0.735000 ;
      RECT 1.915000  1.835000 2.195000 2.635000 ;
      RECT 1.980000  0.085000 2.155000 0.905000 ;
      RECT 2.490000  1.075000 3.500000 1.245000 ;
      RECT 2.490000  1.245000 2.660000 1.445000 ;
      RECT 2.785000  2.135000 3.035000 2.635000 ;
      RECT 2.825000  0.085000 2.995000 0.550000 ;
      RECT 3.625000  1.795000 3.875000 2.635000 ;
      RECT 3.665000  0.085000 3.835000 0.550000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__or2b_4
MACRO sky130_fd_sc_hd__or3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.600000 0.995000 1.425000 1.325000 ;
        RECT 0.600000 1.325000 0.795000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 2.125000 1.275000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.430000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.415000 2.210000 0.760000 ;
        RECT 1.935000 1.495000 2.210000 2.465000 ;
        RECT 2.040000 0.760000 2.210000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.085000 0.310000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.100000  0.305000 0.355000 0.655000 ;
      RECT 0.100000  0.655000 1.765000 0.825000 ;
      RECT 0.105000  1.495000 0.430000 1.785000 ;
      RECT 0.105000  1.785000 1.275000 1.955000 ;
      RECT 0.525000  0.085000 0.855000 0.485000 ;
      RECT 1.025000  0.305000 1.195000 0.655000 ;
      RECT 1.105000  1.495000 1.765000 1.665000 ;
      RECT 1.105000  1.665000 1.275000 1.785000 ;
      RECT 1.365000  0.085000 1.745000 0.485000 ;
      RECT 1.445000  1.835000 1.725000 2.635000 ;
      RECT 1.595000  0.825000 1.765000 0.995000 ;
      RECT 1.595000  0.995000 1.870000 1.325000 ;
      RECT 1.595000  1.325000 1.765000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__or3_1
MACRO sky130_fd_sc_hd__or3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.995000 1.430000 1.325000 ;
        RECT 0.605000 1.325000 0.830000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 2.125000 1.280000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.435000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.940000 0.415000 2.215000 0.760000 ;
        RECT 1.940000 1.495000 2.215000 2.465000 ;
        RECT 2.045000 0.760000 2.215000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.105000  0.305000 0.360000 0.655000 ;
      RECT 0.105000  0.655000 1.770000 0.825000 ;
      RECT 0.105000  1.495000 0.435000 1.785000 ;
      RECT 0.105000  1.785000 1.270000 1.955000 ;
      RECT 0.530000  0.085000 0.860000 0.485000 ;
      RECT 1.030000  0.305000 1.200000 0.655000 ;
      RECT 1.100000  1.495000 1.770000 1.665000 ;
      RECT 1.100000  1.665000 1.270000 1.785000 ;
      RECT 1.370000  0.085000 1.750000 0.485000 ;
      RECT 1.450000  1.835000 1.730000 2.635000 ;
      RECT 1.600000  0.825000 1.770000 0.995000 ;
      RECT 1.600000  0.995000 1.875000 1.325000 ;
      RECT 1.600000  1.325000 1.770000 1.495000 ;
      RECT 2.385000  0.085000 2.675000 0.915000 ;
      RECT 2.385000  1.430000 2.675000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__or3_2
MACRO sky130_fd_sc_hd__or3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225000 1.075000 1.700000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 1.075000 1.055000 1.325000 ;
        RECT 0.595000 1.325000 0.830000 2.050000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.305000 0.265000 2.635000 0.735000 ;
        RECT 2.305000 0.735000 4.055000 0.905000 ;
        RECT 2.345000 1.455000 4.055000 1.625000 ;
        RECT 2.345000 1.625000 2.595000 2.465000 ;
        RECT 3.145000 0.265000 3.475000 0.735000 ;
        RECT 3.185000 1.625000 3.435000 2.465000 ;
        RECT 3.765000 0.905000 4.055000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.255000 0.425000 0.725000 ;
      RECT 0.085000  0.725000 2.090000 0.905000 ;
      RECT 0.085000  1.495000 0.425000 2.295000 ;
      RECT 0.085000  2.295000 1.265000 2.465000 ;
      RECT 0.595000  0.085000 0.765000 0.555000 ;
      RECT 0.935000  0.255000 1.265000 0.725000 ;
      RECT 1.000000  1.495000 2.090000 1.665000 ;
      RECT 1.000000  1.665000 1.265000 2.295000 ;
      RECT 1.435000  0.085000 2.135000 0.555000 ;
      RECT 1.435000  1.835000 2.135000 2.635000 ;
      RECT 1.870000  0.905000 2.090000 1.075000 ;
      RECT 1.870000  1.075000 3.595000 1.245000 ;
      RECT 1.870000  1.245000 2.090000 1.495000 ;
      RECT 2.765000  1.795000 3.015000 2.635000 ;
      RECT 2.805000  0.085000 2.975000 0.555000 ;
      RECT 3.605000  1.795000 3.855000 2.635000 ;
      RECT 3.645000  0.085000 3.815000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__or3_4
MACRO sky130_fd_sc_hd__or3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.995000 2.350000 1.325000 ;
        RECT 1.525000 1.325000 1.770000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585000 2.125000 2.200000 2.455000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.425000 1.325000 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.860000 0.415000 3.135000 0.760000 ;
        RECT 2.860000 1.495000 3.135000 2.465000 ;
        RECT 2.965000 0.760000 3.135000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.905000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 0.515000  0.485000 0.845000 0.905000 ;
      RECT 0.595000  0.905000 0.845000 0.995000 ;
      RECT 0.595000  0.995000 1.310000 1.325000 ;
      RECT 0.595000  1.325000 0.765000 1.885000 ;
      RECT 1.025000  0.255000 1.285000 0.655000 ;
      RECT 1.025000  0.655000 2.690000 0.825000 ;
      RECT 1.025000  1.495000 1.355000 1.785000 ;
      RECT 1.025000  1.785000 2.200000 1.955000 ;
      RECT 1.455000  0.085000 1.785000 0.485000 ;
      RECT 1.955000  0.305000 2.125000 0.655000 ;
      RECT 2.030000  1.495000 2.690000 1.665000 ;
      RECT 2.030000  1.665000 2.200000 1.785000 ;
      RECT 2.295000  0.085000 2.670000 0.485000 ;
      RECT 2.370000  1.835000 2.650000 2.635000 ;
      RECT 2.520000  0.825000 2.690000 0.995000 ;
      RECT 2.520000  0.995000 2.795000 1.325000 ;
      RECT 2.520000  1.325000 2.690000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__or3b_1
MACRO sky130_fd_sc_hd__or3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 1.075000 2.230000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 2.125000 3.135000 2.365000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.640000 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935000 0.265000 1.285000 0.595000 ;
        RECT 0.935000 0.595000 1.105000 1.495000 ;
        RECT 0.935000 1.495000 1.330000 1.700000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.290000 0.345000 0.735000 ;
      RECT 0.085000  0.735000 0.765000 0.905000 ;
      RECT 0.085000  1.810000 0.765000 1.870000 ;
      RECT 0.085000  1.870000 2.660000 1.955000 ;
      RECT 0.085000  1.955000 1.720000 2.040000 ;
      RECT 0.085000  2.040000 0.345000 2.220000 ;
      RECT 0.550000  2.210000 0.910000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.565000 ;
      RECT 0.595000  0.905000 0.765000 1.810000 ;
      RECT 1.275000  0.765000 3.135000 0.825000 ;
      RECT 1.275000  0.825000 2.160000 0.905000 ;
      RECT 1.275000  0.905000 1.595000 0.935000 ;
      RECT 1.275000  0.935000 1.445000 1.325000 ;
      RECT 1.425000  0.735000 3.135000 0.765000 ;
      RECT 1.425000  2.210000 1.755000 2.635000 ;
      RECT 1.520000  0.085000 1.690000 0.565000 ;
      RECT 1.550000  1.785000 2.660000 1.870000 ;
      RECT 1.990000  0.305000 2.160000 0.655000 ;
      RECT 1.990000  0.655000 3.135000 0.735000 ;
      RECT 2.330000  0.085000 2.660000 0.485000 ;
      RECT 2.490000  0.995000 2.790000 1.325000 ;
      RECT 2.490000  1.325000 2.660000 1.785000 ;
      RECT 2.830000  0.305000 3.085000 0.605000 ;
      RECT 2.830000  0.605000 3.135000 0.655000 ;
      RECT 2.830000  1.495000 3.135000 1.925000 ;
      RECT 2.965000  0.825000 3.135000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__or3b_2
MACRO sky130_fd_sc_hd__or3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.400000 1.415000 2.720000 1.700000 ;
        RECT 2.535000 0.995000 2.720000 1.415000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.890000 0.995000 3.200000 1.700000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.640000 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935000 0.735000 2.025000 0.905000 ;
        RECT 0.935000 0.905000 1.105000 1.415000 ;
        RECT 0.935000 1.415000 2.220000 1.700000 ;
        RECT 1.000000 0.285000 1.330000 0.735000 ;
        RECT 1.855000 0.255000 2.090000 0.585000 ;
        RECT 1.855000 0.585000 2.025000 0.735000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.290000 0.345000 0.735000 ;
      RECT 0.085000  0.735000 0.765000 0.905000 ;
      RECT 0.085000  1.810000 0.765000 1.870000 ;
      RECT 0.085000  1.870000 3.620000 2.040000 ;
      RECT 0.085000  2.040000 0.345000 2.220000 ;
      RECT 0.550000  2.210000 0.910000 2.635000 ;
      RECT 0.595000  0.905000 0.765000 1.810000 ;
      RECT 0.620000  0.085000 0.790000 0.565000 ;
      RECT 1.275000  1.075000 2.365000 1.245000 ;
      RECT 1.420000  2.210000 1.750000 2.635000 ;
      RECT 1.500000  0.085000 1.670000 0.565000 ;
      RECT 2.195000  0.720000 4.055000 0.825000 ;
      RECT 2.195000  0.825000 2.400000 0.890000 ;
      RECT 2.195000  0.890000 2.365000 1.075000 ;
      RECT 2.250000  0.655000 4.055000 0.720000 ;
      RECT 2.255000  2.210000 2.595000 2.635000 ;
      RECT 2.260000  0.085000 2.590000 0.485000 ;
      RECT 2.760000  0.305000 2.930000 0.655000 ;
      RECT 3.100000  0.085000 3.490000 0.485000 ;
      RECT 3.390000  0.995000 3.680000 1.325000 ;
      RECT 3.390000  1.325000 3.620000 1.870000 ;
      RECT 3.520000  2.210000 4.055000 2.425000 ;
      RECT 3.660000  0.305000 3.915000 0.605000 ;
      RECT 3.660000  0.605000 4.055000 0.655000 ;
      RECT 3.850000  0.825000 4.055000 2.210000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__or3b_4
MACRO sky130_fd_sc_hd__or4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.490000 0.995000 1.895000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 2.125000 1.745000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 0.995000 1.320000 1.615000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.755000 0.440000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 0.415000 2.675000 0.760000 ;
        RECT 2.405000 1.495000 2.675000 2.465000 ;
        RECT 2.505000 0.760000 2.675000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.090000  1.495000 0.410000 1.785000 ;
      RECT 0.090000  1.785000 1.680000 1.955000 ;
      RECT 0.095000  0.085000 0.425000 0.585000 ;
      RECT 0.625000  0.305000 0.795000 0.655000 ;
      RECT 0.625000  0.655000 2.235000 0.825000 ;
      RECT 0.995000  0.085000 1.325000 0.485000 ;
      RECT 1.495000  0.305000 1.665000 0.655000 ;
      RECT 1.510000  1.495000 2.235000 1.665000 ;
      RECT 1.510000  1.665000 1.680000 1.785000 ;
      RECT 1.835000  0.085000 2.215000 0.485000 ;
      RECT 1.915000  1.835000 2.195000 2.635000 ;
      RECT 2.065000  0.825000 2.235000 0.995000 ;
      RECT 2.065000  0.995000 2.335000 1.325000 ;
      RECT 2.065000  1.325000 2.235000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__or4_1
MACRO sky130_fd_sc_hd__or4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.490000 0.995000 1.895000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 2.125000 1.745000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 0.995000 1.320000 1.615000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.755000 0.440000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 0.415000 2.680000 0.760000 ;
        RECT 2.405000 1.495000 2.680000 2.465000 ;
        RECT 2.510000 0.760000 2.680000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  1.495000 0.410000 1.785000 ;
      RECT 0.085000  1.785000 1.680000 1.955000 ;
      RECT 0.090000  0.085000 0.425000 0.585000 ;
      RECT 0.625000  0.305000 0.795000 0.655000 ;
      RECT 0.625000  0.655000 2.235000 0.825000 ;
      RECT 0.995000  0.085000 1.325000 0.485000 ;
      RECT 1.495000  0.305000 1.665000 0.655000 ;
      RECT 1.510000  1.495000 2.235000 1.665000 ;
      RECT 1.510000  1.665000 1.680000 1.785000 ;
      RECT 1.835000  0.085000 2.215000 0.485000 ;
      RECT 1.915000  1.835000 2.195000 2.635000 ;
      RECT 2.065000  0.825000 2.235000 0.995000 ;
      RECT 2.065000  0.995000 2.340000 1.325000 ;
      RECT 2.065000  1.325000 2.235000 1.495000 ;
      RECT 2.850000  0.085000 3.020000 1.000000 ;
      RECT 2.850000  1.455000 3.020000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__or4_2
MACRO sky130_fd_sc_hd__or4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.840000 0.995000 2.010000 1.445000 ;
        RECT 1.840000 1.445000 2.275000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.280000 0.995000 1.610000 1.450000 ;
        RECT 1.400000 1.450000 1.610000 1.785000 ;
        RECT 1.400000 1.785000 1.720000 2.375000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.880000 0.995000 1.050000 1.620000 ;
        RECT 0.880000 1.620000 1.230000 2.375000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.755000 0.370000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.480000 1.455000 4.055000 1.625000 ;
        RECT 2.480000 1.625000 2.730000 2.465000 ;
        RECT 2.520000 0.255000 2.770000 0.725000 ;
        RECT 2.520000 0.725000 4.055000 0.905000 ;
        RECT 3.280000 0.255000 3.610000 0.725000 ;
        RECT 3.320000 1.625000 3.570000 2.465000 ;
        RECT 3.810000 0.905000 4.055000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.085000 0.310000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.115000  1.495000 0.710000 1.665000 ;
      RECT 0.115000  1.665000 0.450000 2.450000 ;
      RECT 0.120000  0.085000 0.370000 0.585000 ;
      RECT 0.540000  0.655000 2.350000 0.825000 ;
      RECT 0.540000  0.825000 0.710000 1.495000 ;
      RECT 0.700000  0.305000 0.870000 0.655000 ;
      RECT 1.070000  0.085000 1.400000 0.485000 ;
      RECT 1.570000  0.305000 1.740000 0.655000 ;
      RECT 1.960000  0.085000 2.340000 0.485000 ;
      RECT 2.005000  1.795000 2.255000 2.635000 ;
      RECT 2.180000  0.825000 2.350000 1.075000 ;
      RECT 2.180000  1.075000 3.640000 1.245000 ;
      RECT 2.900000  1.795000 3.150000 2.635000 ;
      RECT 2.940000  0.085000 3.110000 0.555000 ;
      RECT 3.740000  1.795000 3.990000 2.635000 ;
      RECT 3.780000  0.085000 3.950000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__or4_4
MACRO sky130_fd_sc_hd__or4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.430000 0.995000 2.810000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 2.125000 2.660000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.520000 0.995000 2.260000 1.615000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.755000 0.425000 1.325000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.320000 0.415000 3.595000 0.760000 ;
        RECT 3.320000 1.495000 3.595000 2.465000 ;
        RECT 3.425000 0.760000 3.595000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.085000 0.425000 0.585000 ;
      RECT 0.085000  1.560000 0.425000 2.635000 ;
      RECT 0.595000  0.305000 0.840000 0.995000 ;
      RECT 0.595000  0.995000 1.250000 1.325000 ;
      RECT 0.595000  1.325000 0.835000 1.920000 ;
      RECT 1.030000  1.495000 1.350000 1.785000 ;
      RECT 1.030000  1.785000 2.660000 1.955000 ;
      RECT 1.035000  0.085000 1.365000 0.585000 ;
      RECT 1.565000  0.305000 1.735000 0.655000 ;
      RECT 1.565000  0.655000 3.150000 0.825000 ;
      RECT 1.910000  0.085000 2.240000 0.485000 ;
      RECT 2.410000  0.305000 2.580000 0.655000 ;
      RECT 2.490000  1.495000 3.150000 1.665000 ;
      RECT 2.490000  1.665000 2.660000 1.785000 ;
      RECT 2.750000  0.085000 3.130000 0.485000 ;
      RECT 2.830000  1.835000 3.110000 2.635000 ;
      RECT 2.980000  0.825000 3.150000 0.995000 ;
      RECT 2.980000  0.995000 3.255000 1.325000 ;
      RECT 2.980000  1.325000 3.150000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__or4b_1
MACRO sky130_fd_sc_hd__or4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.755000 1.075000 2.320000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 2.125000 2.670000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.550000 1.075000 3.550000 1.275000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.435000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935000 0.675000 1.250000 0.680000 ;
        RECT 0.935000 0.680000 1.245000 0.790000 ;
        RECT 0.935000 0.790000 1.105000 1.495000 ;
        RECT 0.935000 1.495000 1.250000 1.825000 ;
        RECT 0.970000 0.260000 1.250000 0.675000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.325000 0.350000 0.735000 ;
      RECT 0.085000  0.735000 0.765000 0.905000 ;
      RECT 0.085000  1.605000 0.765000 1.890000 ;
      RECT 0.510000  1.890000 0.765000 1.995000 ;
      RECT 0.510000  1.995000 1.715000 2.165000 ;
      RECT 0.515000  2.335000 0.845000 2.635000 ;
      RECT 0.595000  0.905000 0.765000 1.605000 ;
      RECT 0.630000  0.085000 0.800000 0.565000 ;
      RECT 1.290000  0.995000 1.585000 1.325000 ;
      RECT 1.415000  0.735000 3.055000 0.905000 ;
      RECT 1.415000  0.905000 1.585000 0.995000 ;
      RECT 1.415000  1.325000 1.585000 1.355000 ;
      RECT 1.415000  1.355000 1.600000 1.370000 ;
      RECT 1.415000  1.370000 1.610000 1.380000 ;
      RECT 1.415000  1.380000 1.620000 1.390000 ;
      RECT 1.415000  1.390000 1.625000 1.400000 ;
      RECT 1.415000  1.400000 1.630000 1.410000 ;
      RECT 1.415000  1.410000 1.645000 1.420000 ;
      RECT 1.415000  1.420000 1.655000 1.425000 ;
      RECT 1.415000  1.425000 1.665000 1.445000 ;
      RECT 1.415000  1.445000 3.560000 1.450000 ;
      RECT 1.420000  1.450000 3.560000 1.615000 ;
      RECT 1.435000  0.085000 1.815000 0.485000 ;
      RECT 1.440000  1.785000 3.030000 1.955000 ;
      RECT 1.440000  1.955000 1.715000 1.995000 ;
      RECT 1.480000  2.335000 1.815000 2.635000 ;
      RECT 1.985000  0.305000 2.155000 0.735000 ;
      RECT 2.385000  0.085000 2.715000 0.485000 ;
      RECT 2.860000  1.955000 3.030000 2.215000 ;
      RECT 2.860000  2.215000 3.345000 2.385000 ;
      RECT 2.885000  0.305000 3.055000 0.735000 ;
      RECT 3.225000  0.085000 3.555000 0.585000 ;
      RECT 3.225000  1.615000 3.560000 1.815000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__or4b_2
MACRO sky130_fd_sc_hd__or4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.755000 0.995000 2.925000 1.445000 ;
        RECT 2.755000 1.445000 3.190000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195000 0.995000 2.525000 1.450000 ;
        RECT 2.335000 1.450000 2.525000 1.785000 ;
        RECT 2.335000 1.785000 2.635000 2.375000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.795000 0.995000 1.965000 1.620000 ;
        RECT 1.795000 1.620000 2.155000 2.375000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.995000 0.445000 1.955000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395000 1.455000 4.965000 1.625000 ;
        RECT 3.395000 1.625000 3.645000 2.465000 ;
        RECT 3.435000 0.255000 3.685000 0.725000 ;
        RECT 3.435000 0.725000 4.965000 0.905000 ;
        RECT 4.195000 0.255000 4.525000 0.725000 ;
        RECT 4.235000 1.625000 4.485000 2.465000 ;
        RECT 4.725000 0.905000 4.965000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.825000 ;
      RECT 0.085000  2.135000 0.365000 2.635000 ;
      RECT 0.595000  0.435000 0.785000 0.905000 ;
      RECT 0.595000  2.065000 0.785000 2.455000 ;
      RECT 0.615000  0.905000 0.785000 0.995000 ;
      RECT 0.615000  0.995000 1.215000 1.325000 ;
      RECT 0.615000  1.325000 0.785000 2.065000 ;
      RECT 1.035000  0.085000 1.285000 0.585000 ;
      RECT 1.035000  1.575000 1.625000 1.745000 ;
      RECT 1.035000  1.745000 1.365000 2.450000 ;
      RECT 1.455000  0.655000 3.265000 0.825000 ;
      RECT 1.455000  0.825000 1.625000 1.575000 ;
      RECT 1.615000  0.305000 1.785000 0.655000 ;
      RECT 1.985000  0.085000 2.315000 0.485000 ;
      RECT 2.485000  0.305000 2.655000 0.655000 ;
      RECT 2.875000  0.085000 3.255000 0.485000 ;
      RECT 2.920000  1.795000 3.170000 2.635000 ;
      RECT 3.095000  0.825000 3.265000 1.075000 ;
      RECT 3.095000  1.075000 4.555000 1.245000 ;
      RECT 3.815000  1.795000 4.065000 2.635000 ;
      RECT 3.855000  0.085000 4.025000 0.555000 ;
      RECT 4.655000  1.795000 4.905000 2.635000 ;
      RECT 4.695000  0.085000 4.865000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__or4b_4
MACRO sky130_fd_sc_hd__or4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615000 0.995000 3.270000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.480000 2.125000 3.120000 2.455000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.695000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.995000 1.235000 1.325000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.780000 0.415000 4.055000 0.760000 ;
        RECT 3.780000 1.495000 4.055000 2.465000 ;
        RECT 3.885000 0.760000 4.055000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.450000 0.400000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.865000 ;
      RECT 0.085000  1.865000 1.915000 2.035000 ;
      RECT 0.085000  2.035000 0.345000 2.455000 ;
      RECT 0.515000  2.205000 0.845000 2.635000 ;
      RECT 0.655000  0.085000 0.825000 0.825000 ;
      RECT 0.990000  1.525000 1.575000 1.695000 ;
      RECT 1.075000  0.450000 1.245000 0.655000 ;
      RECT 1.075000  0.655000 1.575000 0.825000 ;
      RECT 1.405000  0.825000 1.575000 1.075000 ;
      RECT 1.405000  1.075000 1.830000 1.245000 ;
      RECT 1.405000  1.245000 1.575000 1.525000 ;
      RECT 1.470000  0.085000 1.845000 0.485000 ;
      RECT 1.510000  2.205000 2.255000 2.375000 ;
      RECT 1.745000  1.415000 2.395000 1.585000 ;
      RECT 1.745000  1.585000 1.915000 1.865000 ;
      RECT 2.015000  0.305000 2.185000 0.655000 ;
      RECT 2.015000  0.655000 3.610000 0.825000 ;
      RECT 2.085000  1.785000 3.120000 1.955000 ;
      RECT 2.085000  1.955000 2.255000 2.205000 ;
      RECT 2.225000  0.995000 2.395000 1.415000 ;
      RECT 2.370000  0.085000 2.700000 0.485000 ;
      RECT 2.870000  0.305000 3.040000 0.655000 ;
      RECT 2.950000  1.495000 3.610000 1.665000 ;
      RECT 2.950000  1.665000 3.120000 1.785000 ;
      RECT 3.210000  0.085000 3.590000 0.485000 ;
      RECT 3.290000  1.835000 3.570000 2.635000 ;
      RECT 3.440000  0.825000 3.610000 0.995000 ;
      RECT 3.440000  0.995000 3.715000 1.325000 ;
      RECT 3.440000  1.325000 3.610000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__or4bb_1
MACRO sky130_fd_sc_hd__or4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.640000 0.995000 3.295000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 2.125000 3.145000 2.455000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.995000 0.780000 1.695000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.995000 1.240000 1.325000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.415000 4.080000 0.760000 ;
        RECT 3.805000 1.495000 4.080000 2.465000 ;
        RECT 3.910000 0.760000 4.080000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.450000 0.405000 0.825000 ;
      RECT 0.085000  0.825000 0.260000 1.865000 ;
      RECT 0.085000  1.865000 1.940000 2.035000 ;
      RECT 0.085000  2.035000 0.345000 2.455000 ;
      RECT 0.515000  2.205000 0.845000 2.635000 ;
      RECT 0.660000  0.085000 0.830000 0.825000 ;
      RECT 0.995000  1.525000 1.600000 1.695000 ;
      RECT 1.080000  0.450000 1.250000 0.655000 ;
      RECT 1.080000  0.655000 1.600000 0.825000 ;
      RECT 1.410000  0.825000 1.600000 1.075000 ;
      RECT 1.410000  1.075000 1.855000 1.245000 ;
      RECT 1.410000  1.245000 1.600000 1.525000 ;
      RECT 1.495000  0.085000 1.850000 0.485000 ;
      RECT 1.535000  2.205000 2.280000 2.375000 ;
      RECT 1.770000  1.415000 2.420000 1.585000 ;
      RECT 1.770000  1.585000 1.940000 1.865000 ;
      RECT 2.025000  0.305000 2.195000 0.655000 ;
      RECT 2.025000  0.655000 3.635000 0.825000 ;
      RECT 2.110000  1.785000 3.145000 1.955000 ;
      RECT 2.110000  1.955000 2.280000 2.205000 ;
      RECT 2.250000  0.995000 2.420000 1.415000 ;
      RECT 2.395000  0.085000 2.725000 0.485000 ;
      RECT 2.895000  0.305000 3.065000 0.655000 ;
      RECT 2.975000  1.495000 3.635000 1.665000 ;
      RECT 2.975000  1.665000 3.145000 1.785000 ;
      RECT 3.235000  0.085000 3.615000 0.485000 ;
      RECT 3.315000  1.835000 3.595000 2.635000 ;
      RECT 3.465000  0.825000 3.635000 0.995000 ;
      RECT 3.465000  0.995000 3.740000 1.325000 ;
      RECT 3.465000  1.325000 3.635000 1.495000 ;
      RECT 4.250000  0.085000 4.420000 1.025000 ;
      RECT 4.250000  1.440000 4.420000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__or4bb_2
MACRO sky130_fd_sc_hd__or4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.235000 0.995000 3.405000 1.445000 ;
        RECT 3.235000 1.445000 3.670000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.675000 0.995000 3.005000 1.450000 ;
        RECT 2.795000 1.450000 3.005000 1.785000 ;
        RECT 2.795000 1.785000 3.115000 2.375000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.695000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.995000 1.235000 1.325000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.875000 1.455000 5.435000 1.625000 ;
        RECT 3.875000 1.625000 4.125000 2.465000 ;
        RECT 3.915000 0.255000 4.165000 0.725000 ;
        RECT 3.915000 0.725000 5.435000 0.905000 ;
        RECT 4.675000 0.255000 5.005000 0.725000 ;
        RECT 4.715000 1.625000 4.965000 2.465000 ;
        RECT 5.205000 0.905000 5.435000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.450000 0.400000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.865000 ;
      RECT 0.085000  1.865000 1.295000 2.035000 ;
      RECT 0.085000  2.035000 0.345000 2.455000 ;
      RECT 0.515000  2.205000 0.845000 2.635000 ;
      RECT 0.655000  0.085000 0.825000 0.825000 ;
      RECT 0.990000  1.525000 1.595000 1.695000 ;
      RECT 1.075000  0.450000 1.245000 0.655000 ;
      RECT 1.075000  0.655000 1.595000 0.825000 ;
      RECT 1.125000  2.035000 1.295000 2.295000 ;
      RECT 1.125000  2.295000 2.445000 2.465000 ;
      RECT 1.405000  0.825000 1.595000 0.995000 ;
      RECT 1.405000  0.995000 1.695000 1.325000 ;
      RECT 1.405000  1.325000 1.595000 1.525000 ;
      RECT 1.510000  1.955000 2.105000 2.125000 ;
      RECT 1.515000  0.085000 1.845000 0.480000 ;
      RECT 1.935000  0.655000 3.745000 0.825000 ;
      RECT 1.935000  0.825000 2.105000 1.955000 ;
      RECT 2.095000  0.305000 2.265000 0.655000 ;
      RECT 2.275000  0.995000 2.445000 2.295000 ;
      RECT 2.465000  0.085000 2.795000 0.485000 ;
      RECT 2.965000  0.305000 3.135000 0.655000 ;
      RECT 3.355000  0.085000 3.735000 0.485000 ;
      RECT 3.400000  1.795000 3.650000 2.635000 ;
      RECT 3.575000  0.825000 3.745000 1.075000 ;
      RECT 3.575000  1.075000 5.035000 1.245000 ;
      RECT 4.295000  1.795000 4.545000 2.635000 ;
      RECT 4.335000  0.085000 4.505000 0.555000 ;
      RECT 5.135000  1.795000 5.385000 2.635000 ;
      RECT 5.175000  0.085000 5.345000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__or4bb_4
MACRO sky130_fd_sc_hd__probe_p_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__probe_p_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 1.075000 1.240000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1.250000 0.560000 4.270000 2.160000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.095000  1.445000 1.595000 1.615000 ;
      RECT 0.095000  1.615000 0.425000 2.465000 ;
      RECT 0.175000  0.255000 0.345000 0.735000 ;
      RECT 0.175000  0.735000 1.595000 0.905000 ;
      RECT 0.515000  0.085000 0.845000 0.565000 ;
      RECT 0.595000  1.835000 0.765000 2.635000 ;
      RECT 0.935000  1.615000 1.265000 2.465000 ;
      RECT 1.015000  0.260000 1.185000 0.735000 ;
      RECT 1.355000  0.085000 1.685000 0.565000 ;
      RECT 1.420000  0.905000 1.595000 1.075000 ;
      RECT 1.420000  1.075000 4.045000 1.245000 ;
      RECT 1.420000  1.245000 1.595000 1.445000 ;
      RECT 1.435000  1.835000 1.605000 2.635000 ;
      RECT 1.855000  0.255000 2.025000 0.735000 ;
      RECT 1.855000  0.735000 4.545000 0.905000 ;
      RECT 1.855000  1.445000 4.545000 1.615000 ;
      RECT 1.855000  1.615000 2.025000 2.465000 ;
      RECT 2.195000  0.085000 2.525000 0.565000 ;
      RECT 2.195000  1.835000 2.525000 2.635000 ;
      RECT 2.695000  0.255000 2.865000 0.735000 ;
      RECT 2.695000  1.615000 2.865000 2.465000 ;
      RECT 3.035000  0.085000 3.365000 0.565000 ;
      RECT 3.035000  1.835000 3.365000 2.635000 ;
      RECT 3.535000  0.255000 3.705000 0.735000 ;
      RECT 3.535000  1.615000 3.705000 2.465000 ;
      RECT 3.875000  0.085000 4.205000 0.565000 ;
      RECT 3.875000  1.835000 4.205000 2.635000 ;
      RECT 4.290000  0.905000 4.545000 1.055000 ;
      RECT 4.290000  1.055000 4.885000 1.315000 ;
      RECT 4.290000  1.315000 4.545000 1.445000 ;
      RECT 4.375000  0.255000 4.545000 0.735000 ;
      RECT 4.375000  1.615000 4.545000 2.465000 ;
      RECT 4.715000  0.085000 5.045000 0.885000 ;
      RECT 4.715000  1.485000 5.045000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.320000  1.105000 4.490000 1.275000 ;
      RECT 4.680000  1.105000 4.850000 1.275000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
    LAYER met1 ;
      RECT 3.465000 1.060000 4.105000 1.075000 ;
      RECT 3.465000 1.075000 4.910000 1.305000 ;
      RECT 3.465000 1.305000 4.105000 1.320000 ;
    LAYER met2 ;
      RECT 3.445000 1.005000 4.125000 1.375000 ;
    LAYER met3 ;
      RECT 3.395000 1.025000 4.175000 1.355000 ;
    LAYER met4 ;
      RECT 1.370000 0.680000 4.150000 1.860000 ;
    LAYER via ;
      RECT 3.495000 1.060000 3.755000 1.320000 ;
      RECT 3.815000 1.060000 4.075000 1.320000 ;
    LAYER via2 ;
      RECT 3.445000 1.050000 3.725000 1.330000 ;
      RECT 3.845000 1.050000 4.125000 1.330000 ;
    LAYER via3 ;
      RECT 3.425000 1.030000 3.745000 1.350000 ;
      RECT 3.825000 1.030000 4.145000 1.350000 ;
    LAYER via4 ;
      RECT 2.970000 0.680000 4.150000 1.860000 ;
  END
END sky130_fd_sc_hd__probe_p_8
MACRO sky130_fd_sc_hd__probec_p_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__probec_p_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 1.075000 1.240000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT -1.140000 0.770000 0.040000 1.950000 ;
        RECT  1.460000 0.770000 2.640000 1.950000 ;
    END
    PORT
      LAYER met5 ;
        RECT -1.260000  0.560000 2.760000 2.160000 ;
        RECT  1.160000 -1.105000 2.760000 0.560000 ;
        RECT  1.160000  2.160000 2.760000 3.825000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 4.360000 -1.170000 6.675000 0.560000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 4.360000 2.160000 6.675000 3.890000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.095000  1.445000 1.595000 1.615000 ;
      RECT 0.095000  1.615000 0.425000 2.465000 ;
      RECT 0.175000  0.255000 0.345000 0.735000 ;
      RECT 0.175000  0.735000 1.595000 0.905000 ;
      RECT 0.515000  0.085000 0.845000 0.565000 ;
      RECT 0.595000  1.835000 0.765000 2.635000 ;
      RECT 0.935000  1.615000 1.265000 2.465000 ;
      RECT 1.015000  0.260000 1.185000 0.735000 ;
      RECT 1.355000  0.085000 1.685000 0.565000 ;
      RECT 1.420000  0.905000 1.595000 1.075000 ;
      RECT 1.420000  1.075000 4.045000 1.245000 ;
      RECT 1.420000  1.245000 1.595000 1.445000 ;
      RECT 1.435000  1.835000 1.605000 2.635000 ;
      RECT 1.855000  0.255000 2.025000 0.735000 ;
      RECT 1.855000  0.735000 4.545000 0.905000 ;
      RECT 1.855000  1.445000 4.545000 1.615000 ;
      RECT 1.855000  1.615000 2.025000 2.465000 ;
      RECT 2.195000  0.085000 2.525000 0.565000 ;
      RECT 2.195000  1.835000 2.525000 2.635000 ;
      RECT 2.695000  0.255000 2.865000 0.735000 ;
      RECT 2.695000  1.615000 2.865000 2.465000 ;
      RECT 3.035000  0.085000 3.365000 0.565000 ;
      RECT 3.035000  1.835000 3.365000 2.635000 ;
      RECT 3.535000  0.255000 3.705000 0.735000 ;
      RECT 3.535000  1.615000 3.705000 2.465000 ;
      RECT 3.875000  0.085000 4.205000 0.565000 ;
      RECT 3.875000  1.835000 4.205000 2.635000 ;
      RECT 4.290000  0.905000 4.545000 1.055000 ;
      RECT 4.290000  1.055000 4.870000 1.315000 ;
      RECT 4.290000  1.315000 4.545000 1.445000 ;
      RECT 4.375000  0.255000 4.545000 0.735000 ;
      RECT 4.375000  1.615000 4.545000 2.465000 ;
      RECT 4.715000  0.085000 5.045000 0.885000 ;
      RECT 4.715000  1.485000 5.045000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.305000  1.105000 4.475000 1.275000 ;
      RECT 4.665000  1.105000 4.835000 1.275000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 5.520000 -0.130000 ;
      RECT 0.000000 -0.130000 5.840000  0.130000 ;
      RECT 0.000000  0.130000 5.520000  0.240000 ;
      RECT 0.000000  2.480000 5.520000  2.590000 ;
      RECT 0.000000  2.590000 5.840000  2.850000 ;
      RECT 0.000000  2.850000 5.520000  2.960000 ;
      RECT 2.020000  1.060000 2.660000  1.120000 ;
      RECT 2.020000  1.120000 4.895000  1.260000 ;
      RECT 2.020000  1.260000 2.660000  1.320000 ;
      RECT 4.245000  1.075000 4.895000  1.120000 ;
      RECT 4.245000  1.260000 4.895000  1.305000 ;
    LAYER met2 ;
      RECT 1.890000  1.050000 2.660000 1.330000 ;
      RECT 5.135000 -0.140000 5.905000 0.140000 ;
      RECT 5.135000  2.580000 5.905000 2.860000 ;
    LAYER met3 ;
      RECT -0.715000  1.030000 0.065000 1.350000 ;
      RECT  1.885000  1.025000 2.665000 1.355000 ;
      RECT  5.130000 -0.165000 5.910000 0.165000 ;
      RECT  5.130000  2.555000 5.910000 2.885000 ;
    LAYER met4 ;
      RECT 4.930000 -0.895000 6.110000 0.285000 ;
      RECT 4.930000  2.435000 6.110000 3.615000 ;
    LAYER via ;
      RECT 2.050000  1.060000 2.310000 1.320000 ;
      RECT 2.370000  1.060000 2.630000 1.320000 ;
      RECT 5.230000 -0.130000 5.490000 0.130000 ;
      RECT 5.230000  2.590000 5.490000 2.850000 ;
      RECT 5.550000 -0.130000 5.810000 0.130000 ;
      RECT 5.550000  2.590000 5.810000 2.850000 ;
    LAYER via2 ;
      RECT 1.935000  1.050000 2.215000 1.330000 ;
      RECT 2.335000  1.050000 2.615000 1.330000 ;
      RECT 5.180000 -0.140000 5.460000 0.140000 ;
      RECT 5.180000  2.580000 5.460000 2.860000 ;
      RECT 5.580000 -0.140000 5.860000 0.140000 ;
      RECT 5.580000  2.580000 5.860000 2.860000 ;
    LAYER via3 ;
      RECT -0.685000  1.030000 -0.365000 1.350000 ;
      RECT -0.285000  1.030000  0.035000 1.350000 ;
      RECT  1.915000  1.030000  2.235000 1.350000 ;
      RECT  2.315000  1.030000  2.635000 1.350000 ;
      RECT  5.160000 -0.160000  5.480000 0.160000 ;
      RECT  5.160000  2.560000  5.480000 2.880000 ;
      RECT  5.560000 -0.160000  5.880000 0.160000 ;
      RECT  5.560000  2.560000  5.880000 2.880000 ;
  END
END sky130_fd_sc_hd__probec_p_8
MACRO sky130_fd_sc_hd__sdfbbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfbbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.26000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775000 1.405000 4.105000 1.575000 ;
        RECT 3.775000 1.575000 4.060000 1.675000 ;
        RECT 3.825000 1.675000 4.060000 2.375000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.915000 0.255000 14.175000 0.785000 ;
        RECT 13.915000 1.470000 14.175000 2.465000 ;
        RECT 13.965000 0.785000 14.175000 1.470000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.500000 0.255000 12.785000 0.715000 ;
        RECT 12.500000 1.630000 12.785000 2.465000 ;
        RECT 12.605000 0.715000 12.785000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.535000 1.095000 11.990000 1.325000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 1.025000 1.695000 1.685000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.345000 2.155000 0.815000 ;
        RECT 1.935000 0.815000 2.315000 1.150000 ;
        RECT 1.935000 1.150000 2.155000 1.695000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.870000 0.735000 6.295000 0.965000 ;
        RECT 5.870000 0.965000 6.215000 1.065000 ;
      LAYER mcon ;
        RECT 6.125000 0.765000 6.295000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755000 0.735000 10.130000 1.065000 ;
      LAYER mcon ;
        RECT 9.805000 0.765000 9.975000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.065000 0.735000  6.355000 0.780000 ;
        RECT 6.065000 0.780000 10.035000 0.920000 ;
        RECT 6.065000 0.920000  6.355000 0.965000 ;
        RECT 9.745000 0.735000 10.035000 0.780000 ;
        RECT 9.745000 0.920000 10.035000 0.965000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.435000 1.625000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.260000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 14.450000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.260000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.260000 0.085000 ;
      RECT  0.000000  2.635000 14.260000 2.805000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.835000 0.805000 ;
      RECT  0.095000  1.795000  0.835000 1.965000 ;
      RECT  0.095000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.605000  0.805000  0.835000 1.795000 ;
      RECT  1.015000  0.345000  1.235000 2.465000 ;
      RECT  1.430000  0.085000  1.705000 0.635000 ;
      RECT  1.430000  1.885000  1.785000 2.635000 ;
      RECT  2.215000  1.875000  2.575000 2.385000 ;
      RECT  2.325000  0.265000  2.655000 0.595000 ;
      RECT  2.405000  1.295000  3.075000 1.405000 ;
      RECT  2.405000  1.405000  2.670000 1.430000 ;
      RECT  2.405000  1.430000  2.630000 1.465000 ;
      RECT  2.405000  1.465000  2.605000 1.505000 ;
      RECT  2.405000  1.505000  2.575000 1.875000 ;
      RECT  2.460000  1.255000  3.075000 1.295000 ;
      RECT  2.485000  0.595000  2.655000 1.075000 ;
      RECT  2.485000  1.075000  3.075000 1.255000 ;
      RECT  2.760000  1.575000  3.605000 1.745000 ;
      RECT  2.760000  1.745000  3.140000 1.905000 ;
      RECT  2.870000  0.305000  3.040000 0.625000 ;
      RECT  2.870000  0.625000  3.645000 0.765000 ;
      RECT  2.870000  0.765000  3.770000 0.795000 ;
      RECT  2.970000  1.905000  3.140000 2.465000 ;
      RECT  3.225000  0.085000  3.555000 0.445000 ;
      RECT  3.310000  2.215000  3.640000 2.635000 ;
      RECT  3.430000  0.795000  3.770000 1.095000 ;
      RECT  3.430000  1.095000  3.605000 1.575000 ;
      RECT  3.950000  0.425000  4.330000 0.595000 ;
      RECT  3.950000  0.595000  4.120000 1.065000 ;
      RECT  3.950000  1.065000  4.400000 1.105000 ;
      RECT  3.950000  1.105000  4.410000 1.175000 ;
      RECT  3.950000  1.175000  4.445000 1.235000 ;
      RECT  4.160000  0.265000  4.330000 0.425000 ;
      RECT  4.225000  1.235000  4.445000 1.275000 ;
      RECT  4.230000  2.135000  4.445000 2.465000 ;
      RECT  4.245000  1.275000  4.445000 1.305000 ;
      RECT  4.275000  1.305000  4.445000 2.135000 ;
      RECT  4.555000  0.265000  5.655000 0.465000 ;
      RECT  4.570000  0.705000  4.790000 1.035000 ;
      RECT  4.615000  1.035000  4.790000 1.575000 ;
      RECT  4.615000  1.575000  5.125000 1.955000 ;
      RECT  4.635000  2.250000  5.465000 2.420000 ;
      RECT  5.000000  0.735000  5.330000 1.015000 ;
      RECT  5.295000  1.195000  5.670000 1.235000 ;
      RECT  5.295000  1.235000  6.645000 1.405000 ;
      RECT  5.295000  1.405000  5.465000 2.250000 ;
      RECT  5.485000  0.465000  5.655000 0.585000 ;
      RECT  5.485000  0.585000  5.670000 0.655000 ;
      RECT  5.500000  0.655000  5.670000 1.195000 ;
      RECT  5.635000  1.575000  5.885000 1.785000 ;
      RECT  5.635000  1.785000  6.985000 2.035000 ;
      RECT  5.705000  2.205000  6.085000 2.635000 ;
      RECT  5.835000  0.085000  6.005000 0.525000 ;
      RECT  6.260000  0.255000  7.350000 0.425000 ;
      RECT  6.260000  0.425000  6.590000 0.465000 ;
      RECT  6.385000  2.035000  6.555000 2.375000 ;
      RECT  6.395000  1.405000  6.645000 1.485000 ;
      RECT  6.425000  1.155000  6.645000 1.235000 ;
      RECT  6.680000  0.610000  7.010000 0.780000 ;
      RECT  6.810000  0.780000  7.010000 0.895000 ;
      RECT  6.810000  0.895000  8.125000 1.060000 ;
      RECT  6.815000  1.060000  8.125000 1.065000 ;
      RECT  6.815000  1.065000  6.985000 1.785000 ;
      RECT  7.155000  1.235000  7.485000 1.415000 ;
      RECT  7.155000  1.415000  8.160000 1.655000 ;
      RECT  7.175000  1.915000  7.505000 2.635000 ;
      RECT  7.180000  0.425000  7.350000 0.715000 ;
      RECT  7.620000  0.085000  7.975000 0.465000 ;
      RECT  7.795000  1.065000  8.125000 1.235000 ;
      RECT  8.360000  1.575000  8.595000 1.985000 ;
      RECT  8.420000  0.705000  8.705000 1.125000 ;
      RECT  8.420000  1.125000  9.040000 1.305000 ;
      RECT  8.550000  2.250000  9.380000 2.420000 ;
      RECT  8.615000  0.265000  9.380000 0.465000 ;
      RECT  8.835000  1.305000  9.040000 1.905000 ;
      RECT  9.210000  0.465000  9.380000 1.235000 ;
      RECT  9.210000  1.235000 10.560000 1.405000 ;
      RECT  9.210000  1.405000  9.380000 2.250000 ;
      RECT  9.550000  1.575000  9.800000 1.915000 ;
      RECT  9.550000  1.915000 12.330000 2.085000 ;
      RECT  9.560000  0.085000  9.820000 0.525000 ;
      RECT  9.620000  2.255000 10.000000 2.635000 ;
      RECT 10.080000  0.255000 11.250000 0.425000 ;
      RECT 10.080000  0.425000 10.410000 0.545000 ;
      RECT 10.240000  2.085000 10.410000 2.375000 ;
      RECT 10.340000  1.075000 10.560000 1.235000 ;
      RECT 10.575000  0.595000 10.905000 0.780000 ;
      RECT 10.730000  0.780000 10.905000 1.915000 ;
      RECT 10.940000  2.255000 12.330000 2.635000 ;
      RECT 11.075000  0.425000 11.250000 0.585000 ;
      RECT 11.080000  0.755000 11.775000 0.925000 ;
      RECT 11.080000  0.925000 11.355000 1.575000 ;
      RECT 11.080000  1.575000 11.855000 1.745000 ;
      RECT 11.565000  0.265000 11.775000 0.755000 ;
      RECT 12.000000  0.085000 12.330000 0.805000 ;
      RECT 12.160000  0.995000 12.425000 1.325000 ;
      RECT 12.160000  1.325000 12.330000 1.915000 ;
      RECT 12.960000  0.255000 13.275000 0.995000 ;
      RECT 12.960000  0.995000 13.795000 1.325000 ;
      RECT 12.960000  1.325000 13.275000 2.415000 ;
      RECT 13.455000  0.085000 13.745000 0.545000 ;
      RECT 13.455000  1.765000 13.740000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  0.765000  0.775000 0.935000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  1.785000  1.235000 1.955000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  1.105000  3.075000 1.275000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.230000  1.105000  4.400000 1.275000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.785000  4.915000 1.955000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.155000  0.765000  5.325000 0.935000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  1.445000  8.135000 1.615000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  1.105000  8.595000 1.275000 ;
      RECT  8.425000  1.785000  8.595000 1.955000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  1.445000 11.355000 1.615000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
    LAYER met1 ;
      RECT  0.545000 0.735000  0.835000 0.780000 ;
      RECT  0.545000 0.780000  5.385000 0.920000 ;
      RECT  0.545000 0.920000  0.835000 0.965000 ;
      RECT  1.005000 1.755000  1.295000 1.800000 ;
      RECT  1.005000 1.800000  8.655000 1.940000 ;
      RECT  1.005000 1.940000  1.295000 1.985000 ;
      RECT  2.845000 1.075000  3.135000 1.120000 ;
      RECT  2.845000 1.120000  4.460000 1.260000 ;
      RECT  2.845000 1.260000  3.135000 1.305000 ;
      RECT  4.170000 1.075000  4.460000 1.120000 ;
      RECT  4.170000 1.260000  4.460000 1.305000 ;
      RECT  4.685000 1.755000  4.975000 1.800000 ;
      RECT  4.685000 1.940000  4.975000 1.985000 ;
      RECT  5.095000 0.735000  5.385000 0.780000 ;
      RECT  5.095000 0.920000  5.385000 0.965000 ;
      RECT  5.170000 0.965000  5.385000 1.120000 ;
      RECT  5.170000 1.120000  8.655000 1.260000 ;
      RECT  7.905000 1.415000  8.195000 1.460000 ;
      RECT  7.905000 1.460000 11.415000 1.600000 ;
      RECT  7.905000 1.600000  8.195000 1.645000 ;
      RECT  8.365000 1.075000  8.655000 1.120000 ;
      RECT  8.365000 1.260000  8.655000 1.305000 ;
      RECT  8.365000 1.755000  8.655000 1.800000 ;
      RECT  8.365000 1.940000  8.655000 1.985000 ;
      RECT 11.125000 1.415000 11.415000 1.460000 ;
      RECT 11.125000 1.600000 11.415000 1.645000 ;
  END
END sky130_fd_sc_hd__sdfbbn_1
MACRO sky130_fd_sc_hd__sdfbbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfbbn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.18000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825000 1.325000 4.025000 2.375000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.415000 0.255000 14.665000 0.825000 ;
        RECT 14.415000 1.445000 14.665000 2.465000 ;
        RECT 14.460000 0.825000 14.665000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.580000 0.255000 12.830000 0.715000 ;
        RECT 12.580000 1.630000 12.830000 2.465000 ;
        RECT 12.660000 0.715000 12.830000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.590000 1.095000 12.070000 1.325000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 1.025000 1.695000 1.685000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.345000 2.145000 0.765000 ;
        RECT 1.935000 0.765000 2.335000 1.095000 ;
        RECT 1.935000 1.095000 2.155000 1.695000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 0.735000 6.295000 0.965000 ;
        RECT 5.885000 0.965000 6.215000 1.065000 ;
      LAYER mcon ;
        RECT 6.125000 0.765000 6.295000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755000 0.735000 10.130000 1.065000 ;
      LAYER mcon ;
        RECT 9.805000 0.765000 9.975000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.065000 0.735000  6.355000 0.780000 ;
        RECT 6.065000 0.780000 10.035000 0.920000 ;
        RECT 6.065000 0.920000  6.355000 0.965000 ;
        RECT 9.745000 0.735000 10.035000 0.780000 ;
        RECT 9.745000 0.920000 10.035000 0.965000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.435000 1.625000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 15.180000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 15.370000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 15.180000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.180000 0.085000 ;
      RECT  0.000000  2.635000 15.180000 2.805000 ;
      RECT  0.170000  0.345000  0.345000 0.635000 ;
      RECT  0.170000  0.635000  0.835000 0.805000 ;
      RECT  0.170000  1.795000  0.835000 1.965000 ;
      RECT  0.170000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.605000  0.805000  0.835000 1.795000 ;
      RECT  1.015000  0.345000  1.235000 2.465000 ;
      RECT  1.430000  0.085000  1.705000 0.635000 ;
      RECT  1.430000  1.885000  1.785000 2.635000 ;
      RECT  2.215000  1.875000  2.575000 2.385000 ;
      RECT  2.315000  0.265000  2.730000 0.595000 ;
      RECT  2.405000  1.250000  3.075000 1.405000 ;
      RECT  2.405000  1.405000  2.575000 1.875000 ;
      RECT  2.435000  1.235000  3.075000 1.250000 ;
      RECT  2.560000  0.595000  2.730000 1.075000 ;
      RECT  2.560000  1.075000  3.075000 1.235000 ;
      RECT  2.745000  1.575000  3.645000 1.745000 ;
      RECT  2.745000  1.745000  3.065000 1.905000 ;
      RECT  2.895000  1.905000  3.065000 2.465000 ;
      RECT  2.955000  0.305000  3.125000 0.625000 ;
      RECT  2.955000  0.625000  3.645000 0.765000 ;
      RECT  2.955000  0.765000  3.770000 0.795000 ;
      RECT  3.295000  2.215000  3.640000 2.635000 ;
      RECT  3.370000  0.085000  3.700000 0.445000 ;
      RECT  3.475000  0.795000  3.770000 1.095000 ;
      RECT  3.475000  1.095000  3.645000 1.575000 ;
      RECT  4.230000  0.305000  4.455000 2.465000 ;
      RECT  4.625000  0.705000  4.845000 1.575000 ;
      RECT  4.625000  1.575000  5.125000 1.955000 ;
      RECT  4.635000  2.250000  5.465000 2.420000 ;
      RECT  4.700000  0.265000  5.715000 0.465000 ;
      RECT  5.025000  0.645000  5.375000 1.015000 ;
      RECT  5.295000  1.195000  5.715000 1.235000 ;
      RECT  5.295000  1.235000  6.645000 1.405000 ;
      RECT  5.295000  1.405000  5.465000 2.250000 ;
      RECT  5.545000  0.465000  5.715000 1.195000 ;
      RECT  5.635000  1.575000  5.885000 1.785000 ;
      RECT  5.635000  1.785000  6.985000 2.035000 ;
      RECT  5.705000  2.205000  6.085000 2.635000 ;
      RECT  5.885000  0.085000  6.055000 0.525000 ;
      RECT  6.225000  0.255000  7.375000 0.425000 ;
      RECT  6.225000  0.425000  6.555000 0.505000 ;
      RECT  6.385000  2.035000  6.555000 2.375000 ;
      RECT  6.395000  1.405000  6.645000 1.485000 ;
      RECT  6.425000  1.155000  6.645000 1.235000 ;
      RECT  6.705000  0.595000  7.035000 0.765000 ;
      RECT  6.815000  0.765000  7.035000 0.895000 ;
      RECT  6.815000  0.895000  8.125000 1.065000 ;
      RECT  6.815000  1.065000  6.985000 1.785000 ;
      RECT  7.155000  1.235000  7.485000 1.415000 ;
      RECT  7.155000  1.415000  8.160000 1.655000 ;
      RECT  7.175000  1.915000  7.505000 2.635000 ;
      RECT  7.205000  0.425000  7.375000 0.715000 ;
      RECT  7.645000  0.085000  7.975000 0.465000 ;
      RECT  7.795000  1.065000  8.125000 1.235000 ;
      RECT  8.360000  1.575000  8.595000 1.985000 ;
      RECT  8.420000  0.705000  8.705000 1.125000 ;
      RECT  8.420000  1.125000  9.040000 1.305000 ;
      RECT  8.550000  2.250000  9.380000 2.420000 ;
      RECT  8.615000  0.265000  9.380000 0.465000 ;
      RECT  8.835000  1.305000  9.040000 1.905000 ;
      RECT  9.210000  0.465000  9.380000 1.235000 ;
      RECT  9.210000  1.235000 10.560000 1.405000 ;
      RECT  9.210000  1.405000  9.380000 2.250000 ;
      RECT  9.550000  1.575000  9.800000 1.915000 ;
      RECT  9.550000  1.915000 12.410000 2.085000 ;
      RECT  9.560000  0.085000  9.820000 0.525000 ;
      RECT  9.620000  2.255000 10.000000 2.635000 ;
      RECT 10.080000  0.255000 11.250000 0.425000 ;
      RECT 10.080000  0.425000 10.410000 0.545000 ;
      RECT 10.240000  2.085000 10.410000 2.375000 ;
      RECT 10.340000  1.075000 10.560000 1.235000 ;
      RECT 10.580000  0.595000 10.910000 0.780000 ;
      RECT 10.730000  0.780000 10.910000 1.915000 ;
      RECT 10.940000  2.255000 12.410000 2.635000 ;
      RECT 11.080000  0.425000 11.250000 0.585000 ;
      RECT 11.080000  0.755000 11.845000 0.925000 ;
      RECT 11.080000  0.925000 11.355000 1.575000 ;
      RECT 11.080000  1.575000 11.925000 1.745000 ;
      RECT 11.620000  0.265000 11.845000 0.755000 ;
      RECT 12.080000  0.085000 12.410000 0.805000 ;
      RECT 12.240000  0.995000 12.480000 1.325000 ;
      RECT 12.240000  1.325000 12.410000 1.915000 ;
      RECT 13.000000  0.085000 13.235000 0.885000 ;
      RECT 13.000000  1.495000 13.235000 2.635000 ;
      RECT 13.455000  0.255000 13.770000 0.995000 ;
      RECT 13.455000  0.995000 14.290000 1.325000 ;
      RECT 13.455000  1.325000 13.770000 2.415000 ;
      RECT 13.950000  0.085000 14.245000 0.545000 ;
      RECT 13.950000  1.765000 14.245000 2.635000 ;
      RECT 14.835000  0.085000 15.075000 0.885000 ;
      RECT 14.835000  1.495000 15.075000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  0.765000  0.775000 0.935000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  1.785000  1.235000 1.955000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  1.105000  3.075000 1.275000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  1.105000  4.455000 1.275000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.785000  4.915000 1.955000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  0.765000  5.375000 0.935000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  1.445000  8.135000 1.615000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  1.105000  8.595000 1.275000 ;
      RECT  8.425000  1.785000  8.595000 1.955000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  1.445000 11.355000 1.615000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
    LAYER met1 ;
      RECT  0.545000 0.735000  0.835000 0.780000 ;
      RECT  0.545000 0.780000  5.435000 0.920000 ;
      RECT  0.545000 0.920000  0.835000 0.965000 ;
      RECT  1.005000 1.755000  1.295000 1.800000 ;
      RECT  1.005000 1.800000  8.655000 1.940000 ;
      RECT  1.005000 1.940000  1.295000 1.985000 ;
      RECT  2.845000 1.075000  3.135000 1.120000 ;
      RECT  2.845000 1.120000  4.515000 1.260000 ;
      RECT  2.845000 1.260000  3.135000 1.305000 ;
      RECT  4.225000 1.075000  4.515000 1.120000 ;
      RECT  4.225000 1.260000  4.515000 1.305000 ;
      RECT  4.685000 1.755000  4.975000 1.800000 ;
      RECT  4.685000 1.940000  4.975000 1.985000 ;
      RECT  5.145000 0.735000  5.435000 0.780000 ;
      RECT  5.145000 0.920000  5.435000 0.965000 ;
      RECT  5.220000 0.965000  5.435000 1.120000 ;
      RECT  5.220000 1.120000  8.655000 1.260000 ;
      RECT  7.905000 1.415000  8.195000 1.460000 ;
      RECT  7.905000 1.460000 11.415000 1.600000 ;
      RECT  7.905000 1.600000  8.195000 1.645000 ;
      RECT  8.365000 1.075000  8.655000 1.120000 ;
      RECT  8.365000 1.260000  8.655000 1.305000 ;
      RECT  8.365000 1.755000  8.655000 1.800000 ;
      RECT  8.365000 1.940000  8.655000 1.985000 ;
      RECT 11.125000 1.415000 11.415000 1.460000 ;
      RECT 11.125000 1.600000 11.415000 1.645000 ;
  END
END sky130_fd_sc_hd__sdfbbn_2
MACRO sky130_fd_sc_hd__sdfbbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfbbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.26000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825000 1.325000 4.025000 2.375000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.915000 0.255000 14.175000 0.825000 ;
        RECT 13.915000 1.605000 14.175000 2.465000 ;
        RECT 13.965000 0.825000 14.175000 1.605000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.500000 0.255000 12.785000 0.715000 ;
        RECT 12.500000 1.630000 12.785000 2.465000 ;
        RECT 12.605000 0.715000 12.785000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.535000 1.095000 11.990000 1.325000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.440000 1.025000 1.720000 1.685000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.960000 0.345000 2.180000 0.845000 ;
        RECT 1.960000 0.845000 2.415000 1.015000 ;
        RECT 1.960000 1.015000 2.180000 1.695000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 0.735000 6.295000 0.965000 ;
        RECT 5.885000 0.965000 6.215000 1.065000 ;
      LAYER mcon ;
        RECT 6.125000 0.765000 6.295000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755000 0.735000 10.130000 1.065000 ;
      LAYER mcon ;
        RECT 9.805000 0.765000 9.975000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.065000 0.735000  6.355000 0.780000 ;
        RECT 6.065000 0.780000 10.035000 0.920000 ;
        RECT 6.065000 0.920000  6.355000 0.965000 ;
        RECT 9.745000 0.735000 10.035000 0.780000 ;
        RECT 9.745000 0.920000 10.035000 0.965000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.435000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.260000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 14.450000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.260000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.260000 0.085000 ;
      RECT  0.000000  2.635000 14.260000 2.805000 ;
      RECT  0.170000  0.345000  0.345000 0.635000 ;
      RECT  0.170000  0.635000  0.835000 0.805000 ;
      RECT  0.170000  1.795000  0.835000 1.965000 ;
      RECT  0.170000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.605000  0.805000  0.835000 1.795000 ;
      RECT  1.015000  0.345000  1.240000 2.465000 ;
      RECT  1.455000  0.085000  1.705000 0.635000 ;
      RECT  1.455000  1.885000  1.785000 2.635000 ;
      RECT  2.235000  1.875000  2.565000 2.385000 ;
      RECT  2.350000  0.265000  2.755000 0.595000 ;
      RECT  2.350000  1.185000  3.075000 1.365000 ;
      RECT  2.350000  1.365000  2.565000 1.875000 ;
      RECT  2.585000  0.595000  2.755000 1.075000 ;
      RECT  2.585000  1.075000  3.075000 1.185000 ;
      RECT  2.745000  1.575000  3.645000 1.745000 ;
      RECT  2.745000  1.745000  3.065000 1.905000 ;
      RECT  2.895000  1.905000  3.065000 2.465000 ;
      RECT  2.925000  0.305000  3.125000 0.625000 ;
      RECT  2.925000  0.625000  3.645000 0.765000 ;
      RECT  2.925000  0.765000  3.770000 0.795000 ;
      RECT  3.310000  2.215000  3.640000 2.635000 ;
      RECT  3.370000  0.085000  3.700000 0.445000 ;
      RECT  3.475000  0.795000  3.770000 1.095000 ;
      RECT  3.475000  1.095000  3.645000 1.575000 ;
      RECT  4.230000  0.305000  4.455000 2.465000 ;
      RECT  4.625000  0.705000  4.845000 1.575000 ;
      RECT  4.625000  1.575000  5.125000 1.955000 ;
      RECT  4.635000  2.250000  5.465000 2.420000 ;
      RECT  4.700000  0.265000  5.715000 0.465000 ;
      RECT  5.025000  0.645000  5.375000 1.015000 ;
      RECT  5.295000  1.195000  5.715000 1.235000 ;
      RECT  5.295000  1.235000  6.645000 1.405000 ;
      RECT  5.295000  1.405000  5.465000 2.250000 ;
      RECT  5.545000  0.465000  5.715000 1.195000 ;
      RECT  5.635000  1.575000  5.885000 1.785000 ;
      RECT  5.635000  1.785000  6.985000 2.035000 ;
      RECT  5.705000  2.205000  6.085000 2.635000 ;
      RECT  5.885000  0.085000  6.055000 0.525000 ;
      RECT  6.225000  0.255000  7.395000 0.425000 ;
      RECT  6.225000  0.425000  6.555000 0.465000 ;
      RECT  6.385000  2.035000  6.555000 2.375000 ;
      RECT  6.395000  1.405000  6.645000 1.485000 ;
      RECT  6.425000  1.155000  6.645000 1.235000 ;
      RECT  6.700000  0.595000  7.030000 0.765000 ;
      RECT  6.815000  0.765000  7.030000 0.895000 ;
      RECT  6.815000  0.895000  8.125000 1.065000 ;
      RECT  6.815000  1.065000  6.985000 1.785000 ;
      RECT  7.155000  1.235000  7.485000 1.415000 ;
      RECT  7.155000  1.415000  8.160000 1.655000 ;
      RECT  7.175000  1.915000  7.505000 2.635000 ;
      RECT  7.200000  0.425000  7.395000 0.715000 ;
      RECT  7.640000  0.085000  7.975000 0.465000 ;
      RECT  7.795000  1.065000  8.125000 1.235000 ;
      RECT  8.360000  1.575000  8.595000 1.985000 ;
      RECT  8.420000  0.705000  8.705000 1.125000 ;
      RECT  8.420000  1.125000  9.040000 1.305000 ;
      RECT  8.550000  2.250000  9.380000 2.420000 ;
      RECT  8.615000  0.265000  9.380000 0.465000 ;
      RECT  8.835000  1.305000  9.040000 1.905000 ;
      RECT  9.210000  0.465000  9.380000 1.235000 ;
      RECT  9.210000  1.235000 10.560000 1.405000 ;
      RECT  9.210000  1.405000  9.380000 2.250000 ;
      RECT  9.550000  1.575000  9.800000 1.915000 ;
      RECT  9.550000  1.915000 12.330000 2.085000 ;
      RECT  9.560000  0.085000  9.820000 0.525000 ;
      RECT  9.620000  2.255000 10.000000 2.635000 ;
      RECT 10.080000  0.255000 11.250000 0.425000 ;
      RECT 10.080000  0.425000 10.430000 0.465000 ;
      RECT 10.240000  2.085000 10.410000 2.375000 ;
      RECT 10.340000  1.075000 10.560000 1.235000 ;
      RECT 10.575000  0.645000 10.905000 0.815000 ;
      RECT 10.730000  0.815000 10.905000 1.915000 ;
      RECT 10.940000  2.255000 12.330000 2.635000 ;
      RECT 11.075000  0.425000 11.250000 0.585000 ;
      RECT 11.080000  0.755000 11.765000 0.925000 ;
      RECT 11.080000  0.925000 11.355000 1.575000 ;
      RECT 11.080000  1.575000 11.855000 1.745000 ;
      RECT 11.565000  0.265000 11.765000 0.755000 ;
      RECT 12.000000  0.085000 12.330000 0.805000 ;
      RECT 12.160000  0.995000 12.425000 1.325000 ;
      RECT 12.160000  1.325000 12.330000 1.915000 ;
      RECT 12.960000  0.255000 13.275000 0.995000 ;
      RECT 12.960000  0.995000 13.795000 1.325000 ;
      RECT 12.960000  1.325000 13.275000 2.415000 ;
      RECT 13.450000  1.765000 13.745000 2.635000 ;
      RECT 13.455000  0.085000 13.745000 0.545000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  1.785000  0.775000 1.955000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  0.765000  1.235000 0.935000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  1.105000  3.075000 1.275000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  1.105000  4.455000 1.275000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.785000  4.915000 1.955000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  0.765000  5.375000 0.935000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  1.445000  8.135000 1.615000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  1.105000  8.595000 1.275000 ;
      RECT  8.425000  1.785000  8.595000 1.955000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  1.445000 11.355000 1.615000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
    LAYER met1 ;
      RECT  0.545000 1.755000  0.835000 1.800000 ;
      RECT  0.545000 1.800000  8.655000 1.940000 ;
      RECT  0.545000 1.940000  0.835000 1.985000 ;
      RECT  1.005000 0.735000  1.295000 0.780000 ;
      RECT  1.005000 0.780000  5.435000 0.920000 ;
      RECT  1.005000 0.920000  1.295000 0.965000 ;
      RECT  2.845000 1.075000  3.135000 1.120000 ;
      RECT  2.845000 1.120000  4.515000 1.260000 ;
      RECT  2.845000 1.260000  3.135000 1.305000 ;
      RECT  4.225000 1.075000  4.515000 1.120000 ;
      RECT  4.225000 1.260000  4.515000 1.305000 ;
      RECT  4.685000 1.755000  4.975000 1.800000 ;
      RECT  4.685000 1.940000  4.975000 1.985000 ;
      RECT  5.145000 0.735000  5.435000 0.780000 ;
      RECT  5.145000 0.920000  5.435000 0.965000 ;
      RECT  5.220000 0.965000  5.435000 1.120000 ;
      RECT  5.220000 1.120000  8.655000 1.260000 ;
      RECT  7.905000 1.415000  8.195000 1.460000 ;
      RECT  7.905000 1.460000 11.415000 1.600000 ;
      RECT  7.905000 1.600000  8.195000 1.645000 ;
      RECT  8.365000 1.075000  8.655000 1.120000 ;
      RECT  8.365000 1.260000  8.655000 1.305000 ;
      RECT  8.365000 1.755000  8.655000 1.800000 ;
      RECT  8.365000 1.940000  8.655000 1.985000 ;
      RECT 11.125000 1.415000 11.415000 1.460000 ;
      RECT 11.125000 1.600000 11.415000 1.645000 ;
  END
END sky130_fd_sc_hd__sdfbbp_1
MACRO sky130_fd_sc_hd__sdfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.88000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 1.355000 3.120000 1.785000 ;
        RECT 2.865000 1.785000 3.120000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.140000 0.265000 11.400000 0.795000 ;
        RECT 11.140000 1.460000 11.400000 2.325000 ;
        RECT 11.150000 1.445000 11.400000 1.460000 ;
        RECT 11.190000 0.795000 11.400000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.510000 1.560000 12.780000 2.465000 ;
        RECT 12.520000 0.255000 12.780000 0.760000 ;
        RECT 12.600000 0.760000 12.780000 1.560000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505000 0.765000 7.035000 1.045000 ;
      LAYER mcon ;
        RECT 6.865000 0.765000 7.035000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525000 1.065000 10.115000 1.275000 ;
        RECT 9.825000 0.635000 10.115000 1.065000 ;
      LAYER mcon ;
        RECT 9.690000 1.105000  9.860000 1.275000 ;
        RECT 9.945000 0.765000 10.115000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445000 0.735000  7.095000 0.780000 ;
        RECT 6.445000 0.780000 10.175000 0.920000 ;
        RECT 6.445000 0.920000  7.095000 0.965000 ;
        RECT 9.630000 0.920000 10.175000 0.965000 ;
        RECT 9.630000 0.965000  9.920000 1.305000 ;
        RECT 9.885000 0.735000 10.175000 0.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.020000 0.285000 4.275000 0.710000 ;
        RECT 4.020000 0.710000 4.395000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.985000 1.730000 2.465000 ;
        RECT 1.485000 1.070000 1.730000 1.985000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.880000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215000 -0.010000 0.235000 0.015000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  1.970000 1.425000 ;
        RECT -0.190000 1.425000 13.070000 2.910000 ;
        RECT  4.405000 1.305000 13.070000 1.425000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.880000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.880000 0.085000 ;
      RECT  0.000000  2.635000 12.880000 2.805000 ;
      RECT  0.090000  1.795000  0.865000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.835000 0.805000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.530000  2.135000  0.860000 2.635000 ;
      RECT  0.660000  0.805000  0.835000 0.995000 ;
      RECT  0.660000  0.995000  0.975000 1.325000 ;
      RECT  0.660000  1.325000  0.865000 1.795000 ;
      RECT  1.015000  0.345000  1.315000 0.675000 ;
      RECT  1.035000  1.730000  1.315000 1.900000 ;
      RECT  1.035000  1.900000  1.205000 2.465000 ;
      RECT  1.145000  0.675000  1.315000 1.730000 ;
      RECT  1.535000  0.395000  1.705000 0.730000 ;
      RECT  1.535000  0.730000  2.225000 0.900000 ;
      RECT  1.875000  0.085000  2.205000 0.560000 ;
      RECT  1.900000  2.055000  2.150000 2.400000 ;
      RECT  1.980000  1.260000  2.470000 1.455000 ;
      RECT  1.980000  1.455000  2.150000 2.055000 ;
      RECT  2.055000  0.900000  2.225000 0.995000 ;
      RECT  2.055000  0.995000  3.085000 1.185000 ;
      RECT  2.055000  1.185000  2.470000 1.260000 ;
      RECT  2.320000  2.040000  2.490000 2.635000 ;
      RECT  2.395000  0.085000  2.725000 0.825000 ;
      RECT  2.915000  0.255000  3.850000 0.425000 ;
      RECT  2.915000  0.425000  3.085000 0.995000 ;
      RECT  3.255000  0.675000  3.425000 1.015000 ;
      RECT  3.255000  1.015000  3.460000 1.185000 ;
      RECT  3.290000  1.185000  3.460000 1.935000 ;
      RECT  3.290000  1.935000  5.075000 2.105000 ;
      RECT  3.460000  2.105000  3.630000 2.465000 ;
      RECT  3.680000  0.425000  3.850000 1.685000 ;
      RECT  4.300000  2.275000  4.630000 2.635000 ;
      RECT  4.445000  0.085000  4.775000 0.540000 ;
      RECT  4.565000  0.715000  5.145000 0.895000 ;
      RECT  4.565000  0.895000  4.735000 1.935000 ;
      RECT  4.905000  1.065000  5.075000 1.395000 ;
      RECT  4.905000  2.105000  5.075000 2.185000 ;
      RECT  4.905000  2.185000  5.275000 2.435000 ;
      RECT  4.975000  0.335000  5.315000 0.505000 ;
      RECT  4.975000  0.505000  5.145000 0.715000 ;
      RECT  5.245000  1.575000  5.495000 1.955000 ;
      RECT  5.325000  0.705000  5.975000 1.035000 ;
      RECT  5.325000  1.035000  5.495000 1.575000 ;
      RECT  5.470000  2.135000  5.835000 2.465000 ;
      RECT  5.485000  0.305000  6.335000 0.475000 ;
      RECT  5.665000  1.215000  7.375000 1.385000 ;
      RECT  5.665000  1.385000  5.835000 2.135000 ;
      RECT  6.005000  1.935000  7.165000 2.105000 ;
      RECT  6.005000  2.105000  6.175000 2.375000 ;
      RECT  6.165000  0.475000  6.335000 1.215000 ;
      RECT  6.285000  1.595000  7.715000 1.765000 ;
      RECT  6.410000  2.355000  6.740000 2.635000 ;
      RECT  6.915000  0.085000  7.245000 0.545000 ;
      RECT  6.995000  2.105000  7.165000 2.375000 ;
      RECT  7.205000  1.005000  7.375000 1.215000 ;
      RECT  7.375000  2.175000  7.745000 2.635000 ;
      RECT  7.455000  0.275000  7.785000 0.445000 ;
      RECT  7.455000  0.445000  7.715000 0.835000 ;
      RECT  7.455000  1.765000  7.715000 1.835000 ;
      RECT  7.455000  1.835000  8.140000 2.005000 ;
      RECT  7.545000  0.835000  7.715000 1.595000 ;
      RECT  7.885000  0.705000  8.095000 1.495000 ;
      RECT  7.885000  1.495000  8.520000 1.655000 ;
      RECT  7.885000  1.655000  8.870000 1.665000 ;
      RECT  7.970000  2.005000  8.140000 2.465000 ;
      RECT  8.005000  0.255000  8.915000 0.535000 ;
      RECT  8.310000  1.665000  8.870000 1.935000 ;
      RECT  8.310000  1.935000  8.840000 1.955000 ;
      RECT  8.320000  2.125000  9.190000 2.465000 ;
      RECT  8.405000  0.920000  8.575000 1.325000 ;
      RECT  8.745000  0.535000  8.915000 1.315000 ;
      RECT  8.745000  1.315000  9.210000 1.485000 ;
      RECT  9.015000  2.035000  9.210000 2.115000 ;
      RECT  9.015000  2.115000  9.190000 2.125000 ;
      RECT  9.040000  1.485000  9.210000 1.575000 ;
      RECT  9.040000  1.575000 10.205000 1.745000 ;
      RECT  9.040000  1.745000  9.210000 2.035000 ;
      RECT  9.085000  0.085000  9.255000 0.525000 ;
      RECT  9.125000  0.695000  9.655000 0.865000 ;
      RECT  9.125000  0.865000  9.295000 1.145000 ;
      RECT  9.360000  2.195000  9.610000 2.635000 ;
      RECT  9.485000  0.295000 10.515000 0.465000 ;
      RECT  9.485000  0.465000  9.655000 0.695000 ;
      RECT  9.780000  1.915000 10.545000 2.085000 ;
      RECT  9.780000  2.085000  9.950000 2.375000 ;
      RECT 10.120000  2.255000 10.450000 2.635000 ;
      RECT 10.345000  0.465000 10.515000 0.995000 ;
      RECT 10.345000  0.995000 11.020000 1.295000 ;
      RECT 10.375000  1.295000 11.020000 1.325000 ;
      RECT 10.375000  1.325000 10.545000 1.915000 ;
      RECT 10.720000  0.085000 10.890000 0.545000 ;
      RECT 10.720000  1.495000 10.970000 2.635000 ;
      RECT 11.650000  1.535000 12.325000 1.705000 ;
      RECT 11.650000  1.705000 11.830000 2.465000 ;
      RECT 11.660000  0.255000 11.830000 0.635000 ;
      RECT 11.660000  0.635000 12.325000 0.805000 ;
      RECT 12.010000  0.085000 12.340000 0.465000 ;
      RECT 12.010000  1.875000 12.340000 2.635000 ;
      RECT 12.155000  0.805000 12.325000 1.060000 ;
      RECT 12.155000  1.060000 12.430000 1.390000 ;
      RECT 12.155000  1.390000 12.325000 1.535000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.805000  1.105000  0.975000 1.275000 ;
      RECT  1.035000  1.785000  1.205000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.905000  1.105000  5.075000 1.275000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.325000  1.785000  5.495000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.405000  1.105000  8.575000 1.275000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.445000  1.785000  8.615000 1.955000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
    LAYER met1 ;
      RECT 0.745000 1.075000 1.035000 1.120000 ;
      RECT 0.745000 1.120000 8.635000 1.260000 ;
      RECT 0.745000 1.260000 1.035000 1.305000 ;
      RECT 0.970000 1.755000 1.270000 1.800000 ;
      RECT 0.970000 1.800000 8.675000 1.940000 ;
      RECT 0.970000 1.940000 1.270000 1.985000 ;
      RECT 4.845000 1.075000 5.135000 1.120000 ;
      RECT 4.845000 1.260000 5.135000 1.305000 ;
      RECT 5.265000 1.755000 5.555000 1.800000 ;
      RECT 5.265000 1.940000 5.555000 1.985000 ;
      RECT 8.345000 1.075000 8.635000 1.120000 ;
      RECT 8.345000 1.260000 8.635000 1.305000 ;
      RECT 8.385000 1.755000 8.675000 1.800000 ;
      RECT 8.385000 1.940000 8.675000 1.985000 ;
  END
END sky130_fd_sc_hd__sdfrbp_1
MACRO sky130_fd_sc_hd__sdfrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.34000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 1.355000 3.120000 1.785000 ;
        RECT 2.865000 1.785000 3.120000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.575000 0.265000 11.925000 1.695000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.435000 1.535000 12.825000 2.080000 ;
        RECT 12.445000 0.310000 12.825000 0.825000 ;
        RECT 12.525000 2.080000 12.825000 2.465000 ;
        RECT 12.655000 0.825000 12.825000 1.535000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505000 0.765000 7.035000 1.045000 ;
      LAYER mcon ;
        RECT 6.865000 0.765000 7.035000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525000 1.065000 10.115000 1.275000 ;
        RECT 9.825000 0.635000 10.115000 1.065000 ;
      LAYER mcon ;
        RECT 9.690000 1.105000  9.860000 1.275000 ;
        RECT 9.945000 0.765000 10.115000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445000 0.735000  7.095000 0.780000 ;
        RECT 6.445000 0.780000 10.175000 0.920000 ;
        RECT 6.445000 0.920000  7.095000 0.965000 ;
        RECT 9.630000 0.920000 10.175000 0.965000 ;
        RECT 9.630000 0.965000  9.920000 1.305000 ;
        RECT 9.885000 0.735000 10.175000 0.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.020000 0.285000 4.275000 0.710000 ;
        RECT 4.020000 0.710000 4.395000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.985000 1.730000 2.465000 ;
        RECT 1.485000 1.070000 1.730000 1.985000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.340000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215000 -0.010000 0.235000 0.015000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  1.970000 1.425000 ;
        RECT -0.190000 1.425000 13.530000 2.910000 ;
        RECT  4.405000 1.305000 13.530000 1.425000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.340000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.340000 0.085000 ;
      RECT  0.000000  2.635000 13.340000 2.805000 ;
      RECT  0.090000  1.795000  0.865000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.835000 0.805000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.530000  2.135000  0.860000 2.635000 ;
      RECT  0.660000  0.805000  0.835000 0.995000 ;
      RECT  0.660000  0.995000  0.975000 1.325000 ;
      RECT  0.660000  1.325000  0.865000 1.795000 ;
      RECT  1.015000  0.345000  1.315000 0.675000 ;
      RECT  1.035000  1.730000  1.315000 1.900000 ;
      RECT  1.035000  1.900000  1.205000 2.465000 ;
      RECT  1.145000  0.675000  1.315000 1.730000 ;
      RECT  1.535000  0.395000  1.705000 0.730000 ;
      RECT  1.535000  0.730000  2.225000 0.900000 ;
      RECT  1.875000  0.085000  2.205000 0.560000 ;
      RECT  1.900000  2.055000  2.150000 2.400000 ;
      RECT  1.980000  1.260000  2.470000 1.455000 ;
      RECT  1.980000  1.455000  2.150000 2.055000 ;
      RECT  2.055000  0.900000  2.225000 0.995000 ;
      RECT  2.055000  0.995000  3.085000 1.185000 ;
      RECT  2.055000  1.185000  2.470000 1.260000 ;
      RECT  2.320000  2.040000  2.490000 2.635000 ;
      RECT  2.395000  0.085000  2.725000 0.825000 ;
      RECT  2.915000  0.255000  3.850000 0.425000 ;
      RECT  2.915000  0.425000  3.085000 0.995000 ;
      RECT  3.255000  0.675000  3.425000 1.015000 ;
      RECT  3.255000  1.015000  3.460000 1.185000 ;
      RECT  3.290000  1.185000  3.460000 1.935000 ;
      RECT  3.290000  1.935000  5.075000 2.105000 ;
      RECT  3.460000  2.105000  3.630000 2.465000 ;
      RECT  3.680000  0.425000  3.850000 1.685000 ;
      RECT  4.300000  2.275000  4.630000 2.635000 ;
      RECT  4.445000  0.085000  4.775000 0.540000 ;
      RECT  4.565000  0.715000  5.145000 0.895000 ;
      RECT  4.565000  0.895000  4.735000 1.935000 ;
      RECT  4.905000  1.065000  5.075000 1.395000 ;
      RECT  4.905000  2.105000  5.075000 2.185000 ;
      RECT  4.905000  2.185000  5.275000 2.435000 ;
      RECT  4.975000  0.335000  5.315000 0.505000 ;
      RECT  4.975000  0.505000  5.145000 0.715000 ;
      RECT  5.245000  1.575000  5.495000 1.955000 ;
      RECT  5.325000  0.705000  5.975000 1.035000 ;
      RECT  5.325000  1.035000  5.495000 1.575000 ;
      RECT  5.470000  2.135000  5.835000 2.465000 ;
      RECT  5.485000  0.305000  6.335000 0.475000 ;
      RECT  5.665000  1.215000  7.375000 1.385000 ;
      RECT  5.665000  1.385000  5.835000 2.135000 ;
      RECT  6.005000  1.935000  7.165000 2.105000 ;
      RECT  6.005000  2.105000  6.175000 2.375000 ;
      RECT  6.165000  0.475000  6.335000 1.215000 ;
      RECT  6.285000  1.595000  7.715000 1.765000 ;
      RECT  6.410000  2.355000  6.740000 2.635000 ;
      RECT  6.915000  0.085000  7.245000 0.545000 ;
      RECT  6.995000  2.105000  7.165000 2.375000 ;
      RECT  7.205000  1.005000  7.375000 1.215000 ;
      RECT  7.375000  2.175000  7.745000 2.635000 ;
      RECT  7.455000  0.275000  7.785000 0.445000 ;
      RECT  7.455000  0.445000  7.715000 0.835000 ;
      RECT  7.455000  1.765000  7.715000 1.835000 ;
      RECT  7.455000  1.835000  8.140000 2.005000 ;
      RECT  7.545000  0.835000  7.715000 1.595000 ;
      RECT  7.885000  0.705000  8.095000 1.495000 ;
      RECT  7.885000  1.495000  8.520000 1.655000 ;
      RECT  7.885000  1.655000  8.870000 1.665000 ;
      RECT  7.970000  2.005000  8.140000 2.465000 ;
      RECT  8.005000  0.255000  8.915000 0.535000 ;
      RECT  8.310000  1.665000  8.870000 1.935000 ;
      RECT  8.310000  1.935000  8.840000 1.955000 ;
      RECT  8.320000  2.125000  9.190000 2.465000 ;
      RECT  8.405000  0.920000  8.575000 1.325000 ;
      RECT  8.745000  0.535000  8.915000 1.315000 ;
      RECT  8.745000  1.315000  9.210000 1.485000 ;
      RECT  9.015000  2.035000  9.210000 2.115000 ;
      RECT  9.015000  2.115000  9.190000 2.125000 ;
      RECT  9.040000  1.485000  9.210000 1.575000 ;
      RECT  9.040000  1.575000 10.205000 1.745000 ;
      RECT  9.040000  1.745000  9.210000 2.035000 ;
      RECT  9.085000  0.085000  9.255000 0.525000 ;
      RECT  9.125000  0.695000  9.655000 0.865000 ;
      RECT  9.125000  0.865000  9.295000 1.145000 ;
      RECT  9.360000  2.195000  9.610000 2.635000 ;
      RECT  9.485000  0.295000 10.515000 0.465000 ;
      RECT  9.485000  0.465000  9.655000 0.695000 ;
      RECT  9.780000  1.915000 10.545000 2.085000 ;
      RECT  9.780000  2.085000  9.950000 2.375000 ;
      RECT 10.120000  2.255000 10.450000 2.635000 ;
      RECT 10.345000  0.465000 10.515000 1.055000 ;
      RECT 10.345000  1.055000 11.060000 1.295000 ;
      RECT 10.375000  1.295000 11.060000 1.325000 ;
      RECT 10.375000  1.325000 10.545000 1.915000 ;
      RECT 10.715000  0.345000 10.885000 0.715000 ;
      RECT 10.715000  0.715000 11.405000 0.885000 ;
      RECT 10.715000  1.795000 11.405000 1.865000 ;
      RECT 10.715000  1.865000 12.265000 2.035000 ;
      RECT 10.715000  2.035000 10.890000 2.465000 ;
      RECT 11.090000  0.085000 11.365000 0.545000 ;
      RECT 11.090000  2.205000 11.420000 2.635000 ;
      RECT 11.230000  0.885000 11.405000 1.795000 ;
      RECT 11.550000  2.035000 12.265000 2.085000 ;
      RECT 12.025000  2.255000 12.355000 2.635000 ;
      RECT 12.095000  0.995000 12.485000 1.325000 ;
      RECT 12.095000  1.325000 12.265000 1.865000 ;
      RECT 12.105000  0.085000 12.275000 0.825000 ;
      RECT 12.995000  0.085000 13.165000 0.930000 ;
      RECT 12.995000  1.495000 13.245000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.805000  1.105000  0.975000 1.275000 ;
      RECT  1.035000  1.785000  1.205000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.905000  1.105000  5.075000 1.275000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.325000  1.785000  5.495000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.405000  1.105000  8.575000 1.275000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.445000  1.785000  8.615000 1.955000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
    LAYER met1 ;
      RECT 0.745000 1.075000 1.035000 1.120000 ;
      RECT 0.745000 1.120000 8.635000 1.260000 ;
      RECT 0.745000 1.260000 1.035000 1.305000 ;
      RECT 0.970000 1.755000 1.270000 1.800000 ;
      RECT 0.970000 1.800000 8.675000 1.940000 ;
      RECT 0.970000 1.940000 1.270000 1.985000 ;
      RECT 4.845000 1.075000 5.135000 1.120000 ;
      RECT 4.845000 1.260000 5.135000 1.305000 ;
      RECT 5.265000 1.755000 5.555000 1.800000 ;
      RECT 5.265000 1.940000 5.555000 1.985000 ;
      RECT 8.345000 1.075000 8.635000 1.120000 ;
      RECT 8.345000 1.260000 8.635000 1.305000 ;
      RECT 8.385000 1.755000 8.675000 1.800000 ;
      RECT 8.385000 1.940000 8.675000 1.985000 ;
  END
END sky130_fd_sc_hd__sdfrbp_2
MACRO sky130_fd_sc_hd__sdfrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.50000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 1.355000 3.120000 1.785000 ;
        RECT 2.865000 1.785000 3.120000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.140000 0.265000 11.400000 0.795000 ;
        RECT 11.140000 1.460000 11.400000 2.325000 ;
        RECT 11.150000 1.445000 11.400000 1.460000 ;
        RECT 11.190000 0.795000 11.400000 1.445000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505000 0.765000 7.035000 1.045000 ;
      LAYER mcon ;
        RECT 6.865000 0.765000 7.035000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525000 1.065000 10.115000 1.275000 ;
        RECT 9.825000 0.635000 10.115000 1.065000 ;
      LAYER mcon ;
        RECT 9.690000 1.105000  9.860000 1.275000 ;
        RECT 9.945000 0.765000 10.115000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445000 0.735000  7.095000 0.780000 ;
        RECT 6.445000 0.780000 10.175000 0.920000 ;
        RECT 6.445000 0.920000  7.095000 0.965000 ;
        RECT 9.630000 0.920000 10.175000 0.965000 ;
        RECT 9.630000 0.965000  9.920000 1.305000 ;
        RECT 9.885000 0.735000 10.175000 0.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.020000 0.285000 4.275000 0.710000 ;
        RECT 4.020000 0.710000 4.395000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.985000 1.730000 2.465000 ;
        RECT 1.485000 1.070000 1.730000 1.985000 ;
    END
  END SCE
  PIN CLK_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.500000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215000 -0.010000 0.235000 0.015000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  1.970000 1.425000 ;
        RECT -0.190000 1.425000 11.690000 2.910000 ;
        RECT  4.405000 1.305000 11.690000 1.425000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.500000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.500000 0.085000 ;
      RECT  0.000000  2.635000 11.500000 2.805000 ;
      RECT  0.090000  1.795000  0.865000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.835000 0.805000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.530000  2.135000  0.860000 2.635000 ;
      RECT  0.660000  0.805000  0.835000 0.995000 ;
      RECT  0.660000  0.995000  0.975000 1.325000 ;
      RECT  0.660000  1.325000  0.865000 1.795000 ;
      RECT  1.015000  0.345000  1.315000 0.675000 ;
      RECT  1.035000  1.730000  1.315000 1.900000 ;
      RECT  1.035000  1.900000  1.205000 2.465000 ;
      RECT  1.145000  0.675000  1.315000 1.730000 ;
      RECT  1.535000  0.395000  1.705000 0.730000 ;
      RECT  1.535000  0.730000  2.225000 0.900000 ;
      RECT  1.875000  0.085000  2.205000 0.560000 ;
      RECT  1.900000  2.055000  2.150000 2.400000 ;
      RECT  1.980000  1.260000  2.470000 1.455000 ;
      RECT  1.980000  1.455000  2.150000 2.055000 ;
      RECT  2.055000  0.900000  2.225000 0.995000 ;
      RECT  2.055000  0.995000  3.085000 1.185000 ;
      RECT  2.055000  1.185000  2.470000 1.260000 ;
      RECT  2.320000  2.040000  2.490000 2.635000 ;
      RECT  2.395000  0.085000  2.725000 0.825000 ;
      RECT  2.915000  0.255000  3.850000 0.425000 ;
      RECT  2.915000  0.425000  3.085000 0.995000 ;
      RECT  3.255000  0.675000  3.425000 1.015000 ;
      RECT  3.255000  1.015000  3.460000 1.185000 ;
      RECT  3.290000  1.185000  3.460000 1.935000 ;
      RECT  3.290000  1.935000  5.075000 2.105000 ;
      RECT  3.460000  2.105000  3.630000 2.465000 ;
      RECT  3.680000  0.425000  3.850000 1.685000 ;
      RECT  4.300000  2.275000  4.630000 2.635000 ;
      RECT  4.445000  0.085000  4.775000 0.540000 ;
      RECT  4.565000  0.715000  5.145000 0.895000 ;
      RECT  4.565000  0.895000  4.735000 1.935000 ;
      RECT  4.905000  1.065000  5.075000 1.395000 ;
      RECT  4.905000  2.105000  5.075000 2.185000 ;
      RECT  4.905000  2.185000  5.275000 2.435000 ;
      RECT  4.975000  0.335000  5.315000 0.505000 ;
      RECT  4.975000  0.505000  5.145000 0.715000 ;
      RECT  5.245000  1.575000  5.495000 1.955000 ;
      RECT  5.325000  0.705000  5.975000 1.035000 ;
      RECT  5.325000  1.035000  5.495000 1.575000 ;
      RECT  5.470000  2.135000  5.835000 2.465000 ;
      RECT  5.485000  0.305000  6.335000 0.475000 ;
      RECT  5.665000  1.215000  7.375000 1.385000 ;
      RECT  5.665000  1.385000  5.835000 2.135000 ;
      RECT  6.005000  1.935000  7.165000 2.105000 ;
      RECT  6.005000  2.105000  6.175000 2.375000 ;
      RECT  6.165000  0.475000  6.335000 1.215000 ;
      RECT  6.285000  1.595000  7.715000 1.765000 ;
      RECT  6.410000  2.355000  6.740000 2.635000 ;
      RECT  6.915000  0.085000  7.245000 0.545000 ;
      RECT  6.995000  2.105000  7.165000 2.375000 ;
      RECT  7.205000  1.005000  7.375000 1.215000 ;
      RECT  7.375000  2.175000  7.745000 2.635000 ;
      RECT  7.455000  0.275000  7.785000 0.445000 ;
      RECT  7.455000  0.445000  7.715000 0.835000 ;
      RECT  7.455000  1.765000  7.715000 1.835000 ;
      RECT  7.455000  1.835000  8.140000 2.005000 ;
      RECT  7.545000  0.835000  7.715000 1.595000 ;
      RECT  7.885000  0.705000  8.095000 1.495000 ;
      RECT  7.885000  1.495000  8.520000 1.655000 ;
      RECT  7.885000  1.655000  8.870000 1.665000 ;
      RECT  7.970000  2.005000  8.140000 2.465000 ;
      RECT  8.005000  0.255000  8.915000 0.535000 ;
      RECT  8.310000  1.665000  8.870000 1.935000 ;
      RECT  8.310000  1.935000  8.840000 1.955000 ;
      RECT  8.320000  2.125000  9.190000 2.465000 ;
      RECT  8.405000  0.920000  8.575000 1.325000 ;
      RECT  8.745000  0.535000  8.915000 1.315000 ;
      RECT  8.745000  1.315000  9.210000 1.485000 ;
      RECT  9.015000  2.035000  9.210000 2.115000 ;
      RECT  9.015000  2.115000  9.190000 2.125000 ;
      RECT  9.040000  1.485000  9.210000 1.575000 ;
      RECT  9.040000  1.575000 10.205000 1.745000 ;
      RECT  9.040000  1.745000  9.210000 2.035000 ;
      RECT  9.085000  0.085000  9.255000 0.525000 ;
      RECT  9.125000  0.695000  9.655000 0.865000 ;
      RECT  9.125000  0.865000  9.295000 1.145000 ;
      RECT  9.360000  2.195000  9.610000 2.635000 ;
      RECT  9.485000  0.295000 10.515000 0.465000 ;
      RECT  9.485000  0.465000  9.655000 0.695000 ;
      RECT  9.780000  1.915000 10.545000 2.085000 ;
      RECT  9.780000  2.085000  9.950000 2.375000 ;
      RECT 10.120000  2.255000 10.450000 2.635000 ;
      RECT 10.345000  0.465000 10.515000 0.995000 ;
      RECT 10.345000  0.995000 11.020000 1.295000 ;
      RECT 10.375000  1.295000 11.020000 1.325000 ;
      RECT 10.375000  1.325000 10.545000 1.915000 ;
      RECT 10.720000  0.085000 10.890000 0.545000 ;
      RECT 10.720000  1.495000 10.970000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.675000  1.785000  0.845000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.145000  1.105000  1.315000 1.275000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.905000  1.105000  5.075000 1.275000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.325000  1.785000  5.495000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.405000  1.105000  8.575000 1.275000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.445000  1.785000  8.615000 1.955000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
    LAYER met1 ;
      RECT 0.615000 1.755000 0.915000 1.800000 ;
      RECT 0.615000 1.800000 8.675000 1.940000 ;
      RECT 0.615000 1.940000 0.915000 1.985000 ;
      RECT 1.085000 1.075000 1.375000 1.120000 ;
      RECT 1.085000 1.120000 8.635000 1.260000 ;
      RECT 1.085000 1.260000 1.375000 1.305000 ;
      RECT 4.845000 1.075000 5.135000 1.120000 ;
      RECT 4.845000 1.260000 5.135000 1.305000 ;
      RECT 5.265000 1.755000 5.555000 1.800000 ;
      RECT 5.265000 1.940000 5.555000 1.985000 ;
      RECT 8.345000 1.075000 8.635000 1.120000 ;
      RECT 8.345000 1.260000 8.635000 1.305000 ;
      RECT 8.385000 1.755000 8.675000 1.800000 ;
      RECT 8.385000 1.940000 8.675000 1.985000 ;
  END
END sky130_fd_sc_hd__sdfrtn_1
MACRO sky130_fd_sc_hd__sdfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.50000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 1.355000 3.120000 1.785000 ;
        RECT 2.865000 1.785000 3.120000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.140000 0.265000 11.400000 0.795000 ;
        RECT 11.140000 1.460000 11.400000 2.325000 ;
        RECT 11.150000 1.445000 11.400000 1.460000 ;
        RECT 11.190000 0.795000 11.400000 1.445000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505000 0.765000 7.035000 1.045000 ;
      LAYER mcon ;
        RECT 6.865000 0.765000 7.035000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525000 1.065000 10.115000 1.275000 ;
        RECT 9.825000 0.635000 10.115000 1.065000 ;
      LAYER mcon ;
        RECT 9.690000 1.105000  9.860000 1.275000 ;
        RECT 9.945000 0.765000 10.115000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445000 0.735000  7.095000 0.780000 ;
        RECT 6.445000 0.780000 10.175000 0.920000 ;
        RECT 6.445000 0.920000  7.095000 0.965000 ;
        RECT 9.630000 0.920000 10.175000 0.965000 ;
        RECT 9.630000 0.965000  9.920000 1.305000 ;
        RECT 9.885000 0.735000 10.175000 0.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.020000 0.285000 4.275000 0.710000 ;
        RECT 4.020000 0.710000 4.395000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.985000 1.730000 2.465000 ;
        RECT 1.485000 1.070000 1.730000 1.985000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.500000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215000 -0.010000 0.235000 0.015000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  1.970000 1.425000 ;
        RECT -0.190000 1.425000 11.690000 2.910000 ;
        RECT  4.405000 1.305000 11.690000 1.425000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.500000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.500000 0.085000 ;
      RECT  0.000000  2.635000 11.500000 2.805000 ;
      RECT  0.090000  1.795000  0.865000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.835000 0.805000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.530000  2.135000  0.860000 2.635000 ;
      RECT  0.660000  0.805000  0.835000 0.995000 ;
      RECT  0.660000  0.995000  0.975000 1.325000 ;
      RECT  0.660000  1.325000  0.865000 1.795000 ;
      RECT  1.015000  0.345000  1.315000 0.675000 ;
      RECT  1.035000  1.730000  1.315000 1.900000 ;
      RECT  1.035000  1.900000  1.205000 2.465000 ;
      RECT  1.145000  0.675000  1.315000 1.730000 ;
      RECT  1.535000  0.395000  1.705000 0.730000 ;
      RECT  1.535000  0.730000  2.225000 0.900000 ;
      RECT  1.875000  0.085000  2.205000 0.560000 ;
      RECT  1.900000  2.055000  2.150000 2.400000 ;
      RECT  1.980000  1.260000  2.470000 1.455000 ;
      RECT  1.980000  1.455000  2.150000 2.055000 ;
      RECT  2.055000  0.900000  2.225000 0.995000 ;
      RECT  2.055000  0.995000  3.085000 1.185000 ;
      RECT  2.055000  1.185000  2.470000 1.260000 ;
      RECT  2.320000  2.040000  2.490000 2.635000 ;
      RECT  2.395000  0.085000  2.725000 0.825000 ;
      RECT  2.915000  0.255000  3.850000 0.425000 ;
      RECT  2.915000  0.425000  3.085000 0.995000 ;
      RECT  3.255000  0.675000  3.425000 1.015000 ;
      RECT  3.255000  1.015000  3.460000 1.185000 ;
      RECT  3.290000  1.185000  3.460000 1.935000 ;
      RECT  3.290000  1.935000  5.075000 2.105000 ;
      RECT  3.460000  2.105000  3.630000 2.465000 ;
      RECT  3.680000  0.425000  3.850000 1.685000 ;
      RECT  4.300000  2.275000  4.630000 2.635000 ;
      RECT  4.445000  0.085000  4.775000 0.540000 ;
      RECT  4.565000  0.715000  5.145000 0.895000 ;
      RECT  4.565000  0.895000  4.735000 1.935000 ;
      RECT  4.905000  1.065000  5.075000 1.395000 ;
      RECT  4.905000  2.105000  5.075000 2.185000 ;
      RECT  4.905000  2.185000  5.275000 2.435000 ;
      RECT  4.975000  0.335000  5.315000 0.505000 ;
      RECT  4.975000  0.505000  5.145000 0.715000 ;
      RECT  5.245000  1.575000  5.495000 1.955000 ;
      RECT  5.325000  0.705000  5.975000 1.035000 ;
      RECT  5.325000  1.035000  5.495000 1.575000 ;
      RECT  5.470000  2.135000  5.835000 2.465000 ;
      RECT  5.485000  0.305000  6.335000 0.475000 ;
      RECT  5.665000  1.215000  7.375000 1.385000 ;
      RECT  5.665000  1.385000  5.835000 2.135000 ;
      RECT  6.005000  1.935000  7.165000 2.105000 ;
      RECT  6.005000  2.105000  6.175000 2.375000 ;
      RECT  6.165000  0.475000  6.335000 1.215000 ;
      RECT  6.285000  1.595000  7.715000 1.765000 ;
      RECT  6.410000  2.355000  6.740000 2.635000 ;
      RECT  6.915000  0.085000  7.245000 0.545000 ;
      RECT  6.995000  2.105000  7.165000 2.375000 ;
      RECT  7.205000  1.005000  7.375000 1.215000 ;
      RECT  7.375000  2.175000  7.745000 2.635000 ;
      RECT  7.455000  0.275000  7.785000 0.445000 ;
      RECT  7.455000  0.445000  7.715000 0.835000 ;
      RECT  7.455000  1.765000  7.715000 1.835000 ;
      RECT  7.455000  1.835000  8.140000 2.005000 ;
      RECT  7.545000  0.835000  7.715000 1.595000 ;
      RECT  7.885000  0.705000  8.095000 1.495000 ;
      RECT  7.885000  1.495000  8.520000 1.655000 ;
      RECT  7.885000  1.655000  8.870000 1.665000 ;
      RECT  7.970000  2.005000  8.140000 2.465000 ;
      RECT  8.005000  0.255000  8.915000 0.535000 ;
      RECT  8.310000  1.665000  8.870000 1.935000 ;
      RECT  8.310000  1.935000  8.840000 1.955000 ;
      RECT  8.320000  2.125000  9.190000 2.465000 ;
      RECT  8.405000  0.920000  8.575000 1.325000 ;
      RECT  8.745000  0.535000  8.915000 1.315000 ;
      RECT  8.745000  1.315000  9.210000 1.485000 ;
      RECT  9.015000  2.035000  9.210000 2.115000 ;
      RECT  9.015000  2.115000  9.190000 2.125000 ;
      RECT  9.040000  1.485000  9.210000 1.575000 ;
      RECT  9.040000  1.575000 10.205000 1.745000 ;
      RECT  9.040000  1.745000  9.210000 2.035000 ;
      RECT  9.085000  0.085000  9.255000 0.525000 ;
      RECT  9.125000  0.695000  9.655000 0.865000 ;
      RECT  9.125000  0.865000  9.295000 1.145000 ;
      RECT  9.360000  2.195000  9.610000 2.635000 ;
      RECT  9.485000  0.295000 10.515000 0.465000 ;
      RECT  9.485000  0.465000  9.655000 0.695000 ;
      RECT  9.780000  1.915000 10.545000 2.085000 ;
      RECT  9.780000  2.085000  9.950000 2.375000 ;
      RECT 10.120000  2.255000 10.450000 2.635000 ;
      RECT 10.345000  0.465000 10.515000 0.995000 ;
      RECT 10.345000  0.995000 11.020000 1.295000 ;
      RECT 10.375000  1.295000 11.020000 1.325000 ;
      RECT 10.375000  1.325000 10.545000 1.915000 ;
      RECT 10.720000  0.085000 10.890000 0.545000 ;
      RECT 10.720000  1.495000 10.970000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.805000  1.105000  0.975000 1.275000 ;
      RECT  1.035000  1.785000  1.205000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.905000  1.105000  5.075000 1.275000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.325000  1.785000  5.495000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.405000  1.105000  8.575000 1.275000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.445000  1.785000  8.615000 1.955000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
    LAYER met1 ;
      RECT 0.745000 1.075000 1.035000 1.120000 ;
      RECT 0.745000 1.120000 8.635000 1.260000 ;
      RECT 0.745000 1.260000 1.035000 1.305000 ;
      RECT 0.970000 1.755000 1.270000 1.800000 ;
      RECT 0.970000 1.800000 8.675000 1.940000 ;
      RECT 0.970000 1.940000 1.270000 1.985000 ;
      RECT 4.845000 1.075000 5.135000 1.120000 ;
      RECT 4.845000 1.260000 5.135000 1.305000 ;
      RECT 5.265000 1.755000 5.555000 1.800000 ;
      RECT 5.265000 1.940000 5.555000 1.985000 ;
      RECT 8.345000 1.075000 8.635000 1.120000 ;
      RECT 8.345000 1.260000 8.635000 1.305000 ;
      RECT 8.385000 1.755000 8.675000 1.800000 ;
      RECT 8.385000 1.940000 8.675000 1.985000 ;
  END
END sky130_fd_sc_hd__sdfrtp_1
MACRO sky130_fd_sc_hd__sdfrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 1.355000 3.120000 1.785000 ;
        RECT 2.865000 1.785000 3.120000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.140000 0.265000 11.400000 0.795000 ;
        RECT 11.140000 1.460000 11.400000 2.325000 ;
        RECT 11.150000 1.445000 11.400000 1.460000 ;
        RECT 11.190000 0.795000 11.400000 1.445000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505000 0.765000 7.035000 1.045000 ;
      LAYER mcon ;
        RECT 6.865000 0.765000 7.035000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525000 1.065000 10.115000 1.275000 ;
        RECT 9.825000 0.635000 10.115000 1.065000 ;
      LAYER mcon ;
        RECT 9.690000 1.105000  9.860000 1.275000 ;
        RECT 9.945000 0.765000 10.115000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445000 0.735000  7.095000 0.780000 ;
        RECT 6.445000 0.780000 10.175000 0.920000 ;
        RECT 6.445000 0.920000  7.095000 0.965000 ;
        RECT 9.630000 0.920000 10.175000 0.965000 ;
        RECT 9.630000 0.965000  9.920000 1.305000 ;
        RECT 9.885000 0.735000 10.175000 0.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.020000 0.285000 4.275000 0.710000 ;
        RECT 4.020000 0.710000 4.395000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.985000 1.730000 2.465000 ;
        RECT 1.485000 1.070000 1.730000 1.985000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215000 -0.010000 0.235000 0.015000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  1.970000 1.425000 ;
        RECT -0.190000 1.425000 12.150000 2.910000 ;
        RECT  4.405000 1.305000 12.150000 1.425000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.090000  1.795000  0.865000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.835000 0.805000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.530000  2.135000  0.860000 2.635000 ;
      RECT  0.660000  0.805000  0.835000 0.995000 ;
      RECT  0.660000  0.995000  0.975000 1.325000 ;
      RECT  0.660000  1.325000  0.865000 1.795000 ;
      RECT  1.015000  0.345000  1.315000 0.675000 ;
      RECT  1.035000  1.730000  1.315000 1.900000 ;
      RECT  1.035000  1.900000  1.205000 2.465000 ;
      RECT  1.145000  0.675000  1.315000 1.730000 ;
      RECT  1.535000  0.395000  1.705000 0.730000 ;
      RECT  1.535000  0.730000  2.225000 0.900000 ;
      RECT  1.875000  0.085000  2.205000 0.560000 ;
      RECT  1.900000  2.055000  2.150000 2.400000 ;
      RECT  1.980000  1.260000  2.470000 1.455000 ;
      RECT  1.980000  1.455000  2.150000 2.055000 ;
      RECT  2.055000  0.900000  2.225000 0.995000 ;
      RECT  2.055000  0.995000  3.085000 1.185000 ;
      RECT  2.055000  1.185000  2.470000 1.260000 ;
      RECT  2.320000  2.040000  2.490000 2.635000 ;
      RECT  2.395000  0.085000  2.725000 0.825000 ;
      RECT  2.915000  0.255000  3.850000 0.425000 ;
      RECT  2.915000  0.425000  3.085000 0.995000 ;
      RECT  3.255000  0.675000  3.425000 1.015000 ;
      RECT  3.255000  1.015000  3.460000 1.185000 ;
      RECT  3.290000  1.185000  3.460000 1.935000 ;
      RECT  3.290000  1.935000  5.075000 2.105000 ;
      RECT  3.460000  2.105000  3.630000 2.465000 ;
      RECT  3.680000  0.425000  3.850000 1.685000 ;
      RECT  4.300000  2.275000  4.630000 2.635000 ;
      RECT  4.445000  0.085000  4.775000 0.540000 ;
      RECT  4.565000  0.715000  5.145000 0.895000 ;
      RECT  4.565000  0.895000  4.735000 1.935000 ;
      RECT  4.905000  1.065000  5.075000 1.395000 ;
      RECT  4.905000  2.105000  5.075000 2.185000 ;
      RECT  4.905000  2.185000  5.275000 2.435000 ;
      RECT  4.975000  0.335000  5.315000 0.505000 ;
      RECT  4.975000  0.505000  5.145000 0.715000 ;
      RECT  5.245000  1.575000  5.495000 1.955000 ;
      RECT  5.325000  0.705000  5.975000 1.035000 ;
      RECT  5.325000  1.035000  5.495000 1.575000 ;
      RECT  5.470000  2.135000  5.835000 2.465000 ;
      RECT  5.485000  0.305000  6.335000 0.475000 ;
      RECT  5.665000  1.215000  7.375000 1.385000 ;
      RECT  5.665000  1.385000  5.835000 2.135000 ;
      RECT  6.005000  1.935000  7.165000 2.105000 ;
      RECT  6.005000  2.105000  6.175000 2.375000 ;
      RECT  6.165000  0.475000  6.335000 1.215000 ;
      RECT  6.285000  1.595000  7.715000 1.765000 ;
      RECT  6.410000  2.355000  6.740000 2.635000 ;
      RECT  6.915000  0.085000  7.245000 0.545000 ;
      RECT  6.995000  2.105000  7.165000 2.375000 ;
      RECT  7.205000  1.005000  7.375000 1.215000 ;
      RECT  7.375000  2.175000  7.745000 2.635000 ;
      RECT  7.455000  0.275000  7.785000 0.445000 ;
      RECT  7.455000  0.445000  7.715000 0.835000 ;
      RECT  7.455000  1.765000  7.715000 1.835000 ;
      RECT  7.455000  1.835000  8.140000 2.005000 ;
      RECT  7.545000  0.835000  7.715000 1.595000 ;
      RECT  7.885000  0.705000  8.095000 1.495000 ;
      RECT  7.885000  1.495000  8.520000 1.655000 ;
      RECT  7.885000  1.655000  8.870000 1.665000 ;
      RECT  7.970000  2.005000  8.140000 2.465000 ;
      RECT  8.005000  0.255000  8.915000 0.535000 ;
      RECT  8.310000  1.665000  8.870000 1.935000 ;
      RECT  8.310000  1.935000  8.840000 1.955000 ;
      RECT  8.320000  2.125000  9.190000 2.465000 ;
      RECT  8.405000  0.920000  8.575000 1.325000 ;
      RECT  8.745000  0.535000  8.915000 1.315000 ;
      RECT  8.745000  1.315000  9.210000 1.485000 ;
      RECT  9.015000  2.035000  9.210000 2.115000 ;
      RECT  9.015000  2.115000  9.190000 2.125000 ;
      RECT  9.040000  1.485000  9.210000 1.575000 ;
      RECT  9.040000  1.575000 10.205000 1.745000 ;
      RECT  9.040000  1.745000  9.210000 2.035000 ;
      RECT  9.085000  0.085000  9.255000 0.525000 ;
      RECT  9.125000  0.695000  9.655000 0.865000 ;
      RECT  9.125000  0.865000  9.295000 1.145000 ;
      RECT  9.360000  2.195000  9.610000 2.635000 ;
      RECT  9.485000  0.295000 10.515000 0.465000 ;
      RECT  9.485000  0.465000  9.655000 0.695000 ;
      RECT  9.780000  1.915000 10.545000 2.085000 ;
      RECT  9.780000  2.085000  9.950000 2.375000 ;
      RECT 10.120000  2.255000 10.450000 2.635000 ;
      RECT 10.345000  0.465000 10.515000 0.995000 ;
      RECT 10.345000  0.995000 11.020000 1.295000 ;
      RECT 10.375000  1.295000 11.020000 1.325000 ;
      RECT 10.375000  1.325000 10.545000 1.915000 ;
      RECT 10.720000  0.085000 10.890000 0.545000 ;
      RECT 10.720000  1.495000 10.970000 2.635000 ;
      RECT 11.570000  0.085000 11.740000 0.545000 ;
      RECT 11.570000  1.495000 11.820000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.805000  1.105000  0.975000 1.275000 ;
      RECT  1.035000  1.785000  1.205000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.905000  1.105000  5.075000 1.275000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.325000  1.785000  5.495000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.405000  1.105000  8.575000 1.275000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.445000  1.785000  8.615000 1.955000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
    LAYER met1 ;
      RECT 0.745000 1.075000 1.035000 1.120000 ;
      RECT 0.745000 1.120000 8.635000 1.260000 ;
      RECT 0.745000 1.260000 1.035000 1.305000 ;
      RECT 0.970000 1.755000 1.270000 1.800000 ;
      RECT 0.970000 1.800000 8.675000 1.940000 ;
      RECT 0.970000 1.940000 1.270000 1.985000 ;
      RECT 4.845000 1.075000 5.135000 1.120000 ;
      RECT 4.845000 1.260000 5.135000 1.305000 ;
      RECT 5.265000 1.755000 5.555000 1.800000 ;
      RECT 5.265000 1.940000 5.555000 1.985000 ;
      RECT 8.345000 1.075000 8.635000 1.120000 ;
      RECT 8.345000 1.260000 8.635000 1.305000 ;
      RECT 8.385000 1.755000 8.675000 1.800000 ;
      RECT 8.385000 1.940000 8.675000 1.985000 ;
  END
END sky130_fd_sc_hd__sdfrtp_2
MACRO sky130_fd_sc_hd__sdfrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.88000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 1.355000 3.120000 1.785000 ;
        RECT 2.865000 1.785000 3.120000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.140000 0.265000 11.400000 0.795000 ;
        RECT 11.140000 1.460000 11.400000 2.325000 ;
        RECT 11.150000 1.445000 11.400000 1.460000 ;
        RECT 11.190000 0.795000 11.400000 0.995000 ;
        RECT 11.190000 0.995000 12.240000 1.325000 ;
        RECT 11.190000 1.325000 11.400000 1.445000 ;
        RECT 11.990000 0.265000 12.240000 0.995000 ;
        RECT 11.990000 1.325000 12.240000 2.325000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505000 0.765000 7.035000 1.045000 ;
      LAYER mcon ;
        RECT 6.865000 0.765000 7.035000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525000 1.065000 10.115000 1.275000 ;
        RECT 9.825000 0.635000 10.115000 1.065000 ;
      LAYER mcon ;
        RECT 9.690000 1.105000  9.860000 1.275000 ;
        RECT 9.945000 0.765000 10.115000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445000 0.735000  7.095000 0.780000 ;
        RECT 6.445000 0.780000 10.175000 0.920000 ;
        RECT 6.445000 0.920000  7.095000 0.965000 ;
        RECT 9.630000 0.920000 10.175000 0.965000 ;
        RECT 9.630000 0.965000  9.920000 1.305000 ;
        RECT 9.885000 0.735000 10.175000 0.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.020000 0.285000 4.275000 0.710000 ;
        RECT 4.020000 0.710000 4.395000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.985000 1.730000 2.465000 ;
        RECT 1.485000 1.070000 1.730000 1.985000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.880000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215000 -0.010000 0.235000 0.015000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  1.970000 1.425000 ;
        RECT -0.190000 1.425000 13.070000 2.910000 ;
        RECT  4.405000 1.305000 13.070000 1.425000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.880000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.880000 0.085000 ;
      RECT  0.000000  2.635000 12.880000 2.805000 ;
      RECT  0.090000  1.795000  0.865000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.835000 0.805000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.530000  2.135000  0.860000 2.635000 ;
      RECT  0.660000  0.805000  0.835000 0.995000 ;
      RECT  0.660000  0.995000  0.975000 1.325000 ;
      RECT  0.660000  1.325000  0.865000 1.795000 ;
      RECT  1.015000  0.345000  1.315000 0.675000 ;
      RECT  1.035000  1.730000  1.315000 1.900000 ;
      RECT  1.035000  1.900000  1.205000 2.465000 ;
      RECT  1.145000  0.675000  1.315000 1.730000 ;
      RECT  1.535000  0.395000  1.705000 0.730000 ;
      RECT  1.535000  0.730000  2.225000 0.900000 ;
      RECT  1.875000  0.085000  2.205000 0.560000 ;
      RECT  1.900000  2.055000  2.150000 2.400000 ;
      RECT  1.980000  1.260000  2.470000 1.455000 ;
      RECT  1.980000  1.455000  2.150000 2.055000 ;
      RECT  2.055000  0.900000  2.225000 0.995000 ;
      RECT  2.055000  0.995000  3.085000 1.185000 ;
      RECT  2.055000  1.185000  2.470000 1.260000 ;
      RECT  2.320000  2.040000  2.490000 2.635000 ;
      RECT  2.395000  0.085000  2.725000 0.825000 ;
      RECT  2.915000  0.255000  3.850000 0.425000 ;
      RECT  2.915000  0.425000  3.085000 0.995000 ;
      RECT  3.255000  0.675000  3.425000 1.015000 ;
      RECT  3.255000  1.015000  3.460000 1.185000 ;
      RECT  3.290000  1.185000  3.460000 1.935000 ;
      RECT  3.290000  1.935000  5.075000 2.105000 ;
      RECT  3.460000  2.105000  3.630000 2.465000 ;
      RECT  3.680000  0.425000  3.850000 1.685000 ;
      RECT  4.300000  2.275000  4.630000 2.635000 ;
      RECT  4.445000  0.085000  4.775000 0.540000 ;
      RECT  4.565000  0.715000  5.145000 0.895000 ;
      RECT  4.565000  0.895000  4.735000 1.935000 ;
      RECT  4.905000  1.065000  5.075000 1.395000 ;
      RECT  4.905000  2.105000  5.075000 2.185000 ;
      RECT  4.905000  2.185000  5.275000 2.435000 ;
      RECT  4.975000  0.335000  5.315000 0.505000 ;
      RECT  4.975000  0.505000  5.145000 0.715000 ;
      RECT  5.245000  1.575000  5.495000 1.955000 ;
      RECT  5.325000  0.705000  5.975000 1.035000 ;
      RECT  5.325000  1.035000  5.495000 1.575000 ;
      RECT  5.470000  2.135000  5.835000 2.465000 ;
      RECT  5.485000  0.305000  6.335000 0.475000 ;
      RECT  5.665000  1.215000  7.375000 1.385000 ;
      RECT  5.665000  1.385000  5.835000 2.135000 ;
      RECT  6.005000  1.935000  7.165000 2.105000 ;
      RECT  6.005000  2.105000  6.175000 2.375000 ;
      RECT  6.165000  0.475000  6.335000 1.215000 ;
      RECT  6.285000  1.595000  7.715000 1.765000 ;
      RECT  6.410000  2.355000  6.740000 2.635000 ;
      RECT  6.915000  0.085000  7.245000 0.545000 ;
      RECT  6.995000  2.105000  7.165000 2.375000 ;
      RECT  7.205000  1.005000  7.375000 1.215000 ;
      RECT  7.375000  2.175000  7.745000 2.635000 ;
      RECT  7.455000  0.275000  7.785000 0.445000 ;
      RECT  7.455000  0.445000  7.715000 0.835000 ;
      RECT  7.455000  1.765000  7.715000 1.835000 ;
      RECT  7.455000  1.835000  8.140000 2.005000 ;
      RECT  7.545000  0.835000  7.715000 1.595000 ;
      RECT  7.885000  0.705000  8.095000 1.495000 ;
      RECT  7.885000  1.495000  8.520000 1.655000 ;
      RECT  7.885000  1.655000  8.870000 1.665000 ;
      RECT  7.970000  2.005000  8.140000 2.465000 ;
      RECT  8.005000  0.255000  8.915000 0.535000 ;
      RECT  8.310000  1.665000  8.870000 1.935000 ;
      RECT  8.310000  1.935000  8.840000 1.955000 ;
      RECT  8.320000  2.125000  9.190000 2.465000 ;
      RECT  8.405000  0.920000  8.575000 1.325000 ;
      RECT  8.745000  0.535000  8.915000 1.315000 ;
      RECT  8.745000  1.315000  9.210000 1.485000 ;
      RECT  9.015000  2.035000  9.210000 2.115000 ;
      RECT  9.015000  2.115000  9.190000 2.125000 ;
      RECT  9.040000  1.485000  9.210000 1.575000 ;
      RECT  9.040000  1.575000 10.205000 1.745000 ;
      RECT  9.040000  1.745000  9.210000 2.035000 ;
      RECT  9.085000  0.085000  9.255000 0.525000 ;
      RECT  9.125000  0.695000  9.655000 0.865000 ;
      RECT  9.125000  0.865000  9.295000 1.145000 ;
      RECT  9.360000  2.195000  9.610000 2.635000 ;
      RECT  9.485000  0.295000 10.515000 0.465000 ;
      RECT  9.485000  0.465000  9.655000 0.695000 ;
      RECT  9.780000  1.915000 10.545000 2.085000 ;
      RECT  9.780000  2.085000  9.950000 2.375000 ;
      RECT 10.120000  2.255000 10.450000 2.635000 ;
      RECT 10.345000  0.465000 10.515000 0.995000 ;
      RECT 10.345000  0.995000 11.020000 1.295000 ;
      RECT 10.375000  1.295000 11.020000 1.325000 ;
      RECT 10.375000  1.325000 10.545000 1.915000 ;
      RECT 10.720000  0.085000 10.890000 0.545000 ;
      RECT 10.720000  1.495000 10.970000 2.635000 ;
      RECT 11.570000  0.085000 11.740000 0.545000 ;
      RECT 11.570000  1.495000 11.820000 2.635000 ;
      RECT 12.410000  0.085000 12.580000 0.545000 ;
      RECT 12.410000  1.495000 12.660000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.805000  1.105000  0.975000 1.275000 ;
      RECT  1.035000  1.785000  1.205000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.905000  1.105000  5.075000 1.275000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.325000  1.785000  5.495000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.405000  1.105000  8.575000 1.275000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.445000  1.785000  8.615000 1.955000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
    LAYER met1 ;
      RECT 0.745000 1.075000 1.035000 1.120000 ;
      RECT 0.745000 1.120000 8.635000 1.260000 ;
      RECT 0.745000 1.260000 1.035000 1.305000 ;
      RECT 0.970000 1.755000 1.270000 1.800000 ;
      RECT 0.970000 1.800000 8.675000 1.940000 ;
      RECT 0.970000 1.940000 1.270000 1.985000 ;
      RECT 4.845000 1.075000 5.135000 1.120000 ;
      RECT 4.845000 1.260000 5.135000 1.305000 ;
      RECT 5.265000 1.755000 5.555000 1.800000 ;
      RECT 5.265000 1.940000 5.555000 1.985000 ;
      RECT 8.345000 1.075000 8.635000 1.120000 ;
      RECT 8.345000 1.260000 8.635000 1.305000 ;
      RECT 8.385000 1.755000 8.675000 1.800000 ;
      RECT 8.385000 1.940000 8.675000 1.985000 ;
  END
END sky130_fd_sc_hd__sdfrtp_4
MACRO sky130_fd_sc_hd__sdfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfsbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.34000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 0.765000 1.335000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.915000 0.275000 13.255000 0.825000 ;
        RECT 12.915000 1.495000 13.255000 2.450000 ;
        RECT 13.070000 0.825000 13.255000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.500000 0.255000 11.830000 2.465000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.345000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.765000 0.825000 1.675000 ;
      LAYER mcon ;
        RECT 0.610000 1.105000 0.780000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.370000 1.075000 2.700000 1.600000 ;
      LAYER mcon ;
        RECT 2.445000 1.105000 2.615000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.550000 1.075000 0.840000 1.120000 ;
        RECT 0.550000 1.120000 2.675000 1.260000 ;
        RECT 0.550000 1.260000 0.840000 1.305000 ;
        RECT 2.385000 1.075000 2.675000 1.120000 ;
        RECT 2.385000 1.260000 2.675000 1.305000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 1.445000 7.015000 1.765000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.885000 1.415000  9.110000 1.525000 ;
        RECT 8.885000 1.525000 10.075000 1.725000 ;
      LAYER mcon ;
        RECT 8.885000 1.445000 9.055000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.580000 1.415000 6.870000 1.460000 ;
        RECT 6.580000 1.460000 9.115000 1.600000 ;
        RECT 6.580000 1.600000 6.870000 1.645000 ;
        RECT 8.825000 1.415000 9.115000 1.460000 ;
        RECT 8.825000 1.600000 9.115000 1.645000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.725000 3.100000 1.055000 ;
        RECT 2.905000 1.055000 3.565000 1.590000 ;
        RECT 2.905000 1.590000 3.085000 1.960000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.340000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 13.530000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.340000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.340000 0.085000 ;
      RECT  0.000000  2.635000 13.340000 2.805000 ;
      RECT  0.085000  0.085000  0.480000 0.595000 ;
      RECT  0.085000  1.845000  1.105000 2.025000 ;
      RECT  0.085000  2.025000  0.345000 2.465000 ;
      RECT  0.515000  2.195000  0.765000 2.635000 ;
      RECT  0.875000  0.280000  1.655000 0.560000 ;
      RECT  0.935000  2.025000  1.105000 2.255000 ;
      RECT  0.935000  2.255000  2.045000 2.465000 ;
      RECT  1.295000  1.870000  1.695000 2.075000 ;
      RECT  1.380000  0.560000  1.655000 0.590000 ;
      RECT  1.380000  0.590000  1.660000 0.600000 ;
      RECT  1.395000  0.600000  1.660000 0.605000 ;
      RECT  1.405000  0.605000  1.660000 0.610000 ;
      RECT  1.420000  0.610000  1.660000 0.615000 ;
      RECT  1.430000  0.615000  1.670000 0.620000 ;
      RECT  1.440000  0.620000  1.670000 0.630000 ;
      RECT  1.445000  0.630000  1.670000 0.635000 ;
      RECT  1.460000  0.635000  1.670000 0.645000 ;
      RECT  1.475000  0.645000  1.670000 0.655000 ;
      RECT  1.475000  0.655000  1.695000 0.665000 ;
      RECT  1.495000  0.665000  1.695000 0.705000 ;
      RECT  1.505000  0.705000  1.695000 1.870000 ;
      RECT  1.825000  0.085000  2.005000 0.545000 ;
      RECT  1.865000  0.715000  2.515000 0.905000 ;
      RECT  1.865000  0.905000  2.200000 1.770000 ;
      RECT  1.865000  1.770000  2.520000 2.085000 ;
      RECT  2.260000  0.255000  2.515000 0.715000 ;
      RECT  2.270000  2.085000  2.520000 2.465000 ;
      RECT  2.690000  0.085000  3.030000 0.555000 ;
      RECT  2.690000  2.140000  3.030000 2.635000 ;
      RECT  3.255000  1.775000  3.995000 1.955000 ;
      RECT  3.255000  1.955000  3.425000 2.325000 ;
      RECT  3.270000  0.255000  3.455000 0.715000 ;
      RECT  3.270000  0.715000  3.995000 0.885000 ;
      RECT  3.595000  2.275000  3.925000 2.635000 ;
      RECT  3.630000  0.085000  3.940000 0.545000 ;
      RECT  3.735000  0.885000  3.995000 1.775000 ;
      RECT  4.095000  2.135000  4.440000 2.465000 ;
      RECT  4.110000  0.255000  4.335000 0.585000 ;
      RECT  4.165000  0.585000  4.335000 1.090000 ;
      RECT  4.165000  1.090000  4.490000 1.420000 ;
      RECT  4.165000  1.420000  4.440000 2.135000 ;
      RECT  4.505000  0.255000  4.830000 0.920000 ;
      RECT  4.610000  1.590000  4.915000 1.615000 ;
      RECT  4.610000  1.615000  4.830000 2.465000 ;
      RECT  4.660000  0.920000  4.830000 1.445000 ;
      RECT  4.660000  1.445000  4.915000 1.590000 ;
      RECT  5.000000  0.255000  5.440000 1.225000 ;
      RECT  5.000000  1.225000  7.660000 1.275000 ;
      RECT  5.030000  2.135000  5.755000 2.465000 ;
      RECT  5.085000  1.275000  6.435000 1.395000 ;
      RECT  5.205000  1.575000  5.415000 1.955000 ;
      RECT  5.585000  1.395000  5.755000 2.135000 ;
      RECT  5.610000  0.085000  6.095000 0.465000 ;
      RECT  5.610000  0.635000  6.535000 0.805000 ;
      RECT  5.610000  0.805000  5.975000 1.015000 ;
      RECT  5.925000  1.575000  6.095000 1.935000 ;
      RECT  5.925000  1.935000  6.765000 2.105000 ;
      RECT  5.945000  2.275000  6.275000 2.635000 ;
      RECT  6.250000  0.975000  7.660000 1.225000 ;
      RECT  6.275000  0.255000  6.535000 0.635000 ;
      RECT  6.550000  2.105000  6.765000 2.450000 ;
      RECT  6.735000  0.085000  7.630000 0.805000 ;
      RECT  7.005000  2.125000  7.960000 2.635000 ;
      RECT  7.190000  1.495000  8.005000 1.955000 ;
      RECT  7.300000  1.275000  7.660000 1.325000 ;
      RECT  7.835000  0.695000  9.040000 0.895000 ;
      RECT  7.835000  0.895000  8.005000 1.495000 ;
      RECT  8.130000  2.125000  8.935000 2.460000 ;
      RECT  8.365000  1.075000  8.595000 1.905000 ;
      RECT  8.410000  0.275000  9.825000 0.445000 ;
      RECT  8.765000  1.895000 10.465000 2.065000 ;
      RECT  8.765000  2.065000  8.935000 2.125000 ;
      RECT  8.810000  0.895000  9.040000 1.245000 ;
      RECT  9.195000  2.235000  9.525000 2.635000 ;
      RECT  9.290000  0.855000  9.465000 1.185000 ;
      RECT  9.290000  1.185000 10.895000 1.355000 ;
      RECT  9.655000  0.445000  9.825000 0.845000 ;
      RECT  9.655000  0.845000 10.545000 1.015000 ;
      RECT  9.695000  2.065000  9.910000 2.450000 ;
      RECT 10.135000  2.235000 10.465000 2.635000 ;
      RECT 10.220000  0.085000 10.390000 0.545000 ;
      RECT 10.245000  1.525000 10.465000 1.895000 ;
      RECT 10.560000  0.255000 10.895000 0.540000 ;
      RECT 10.635000  1.355000 10.895000 2.465000 ;
      RECT 10.715000  0.540000 10.895000 1.185000 ;
      RECT 11.120000  0.085000 11.330000 0.885000 ;
      RECT 11.120000  1.485000 11.330000 2.635000 ;
      RECT 12.060000  0.255000 12.270000 0.995000 ;
      RECT 12.060000  0.995000 12.900000 1.325000 ;
      RECT 12.060000  1.325000 12.270000 2.465000 ;
      RECT 12.540000  0.085000 12.745000 0.825000 ;
      RECT 12.575000  1.575000 12.745000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  1.445000  1.695000 1.615000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  1.785000  3.995000 1.955000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  1.105000  4.455000 1.275000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.445000  4.915000 1.615000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  1.785000  7.675000 1.955000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  1.105000  8.595000 1.275000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
    LAYER met1 ;
      RECT 1.465000 1.415000 1.755000 1.460000 ;
      RECT 1.465000 1.460000 4.975000 1.600000 ;
      RECT 1.465000 1.600000 1.755000 1.645000 ;
      RECT 3.765000 1.755000 4.055000 1.800000 ;
      RECT 3.765000 1.800000 7.735000 1.940000 ;
      RECT 3.765000 1.940000 4.055000 1.985000 ;
      RECT 4.225000 1.075000 4.515000 1.120000 ;
      RECT 4.225000 1.120000 8.655000 1.260000 ;
      RECT 4.225000 1.260000 4.515000 1.305000 ;
      RECT 4.685000 1.415000 4.975000 1.460000 ;
      RECT 4.685000 1.600000 4.975000 1.645000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 7.445000 1.755000 7.735000 1.800000 ;
      RECT 7.445000 1.940000 7.735000 1.985000 ;
      RECT 8.365000 1.075000 8.655000 1.120000 ;
      RECT 8.365000 1.260000 8.655000 1.305000 ;
  END
END sky130_fd_sc_hd__sdfsbp_1
MACRO sky130_fd_sc_hd__sdfsbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfsbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.26000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.765000 1.335000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.410000 0.275000 13.740000 0.825000 ;
        RECT 13.410000 1.495000 13.740000 2.450000 ;
        RECT 13.515000 0.825000 13.740000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.460000 0.255000 11.855000 2.465000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.340000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 0.765000 0.820000 1.675000 ;
      LAYER mcon ;
        RECT 0.605000 1.105000 0.775000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.405000 1.075000 2.735000 1.590000 ;
      LAYER mcon ;
        RECT 2.445000 1.105000 2.615000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.545000 1.075000 0.835000 1.120000 ;
        RECT 0.545000 1.120000 2.675000 1.260000 ;
        RECT 0.545000 1.260000 0.835000 1.305000 ;
        RECT 2.385000 1.075000 2.675000 1.120000 ;
        RECT 2.385000 1.260000 2.675000 1.305000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 1.445000 7.065000 1.765000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.880000 1.435000 9.115000 1.525000 ;
        RECT 8.880000 1.525000 9.935000 1.725000 ;
      LAYER mcon ;
        RECT 8.940000 1.445000 9.110000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.580000 1.415000 6.870000 1.460000 ;
        RECT 6.580000 1.460000 9.170000 1.600000 ;
        RECT 6.580000 1.600000 6.870000 1.645000 ;
        RECT 8.880000 1.415000 9.170000 1.460000 ;
        RECT 8.880000 1.600000 9.170000 1.645000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.725000 3.100000 1.055000 ;
        RECT 2.905000 1.055000 3.565000 1.615000 ;
        RECT 2.905000 1.615000 3.100000 1.970000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.260000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 14.450000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.260000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.260000 0.085000 ;
      RECT  0.000000  2.635000 14.260000 2.805000 ;
      RECT  0.085000  0.085000  0.700000 0.595000 ;
      RECT  0.085000  1.845000  1.185000 2.075000 ;
      RECT  0.085000  2.075000  0.345000 2.465000 ;
      RECT  0.515000  2.275000  0.845000 2.635000 ;
      RECT  0.870000  0.255000  1.670000 0.595000 ;
      RECT  1.015000  2.075000  1.185000 2.255000 ;
      RECT  1.015000  2.255000  2.105000 2.465000 ;
      RECT  1.355000  1.845000  1.695000 2.085000 ;
      RECT  1.495000  0.595000  1.670000 0.645000 ;
      RECT  1.495000  0.645000  1.695000 0.705000 ;
      RECT  1.500000  0.705000  1.695000 0.720000 ;
      RECT  1.505000  0.720000  1.695000 1.845000 ;
      RECT  1.840000  0.085000  2.090000 0.545000 ;
      RECT  1.980000  0.715000  2.530000 0.905000 ;
      RECT  1.980000  0.905000  2.235000 1.760000 ;
      RECT  1.980000  1.760000  2.535000 2.085000 ;
      RECT  2.260000  0.255000  2.530000 0.715000 ;
      RECT  2.275000  2.085000  2.535000 2.465000 ;
      RECT  2.700000  0.085000  3.100000 0.555000 ;
      RECT  2.705000  2.140000  3.100000 2.635000 ;
      RECT  3.270000  0.255000  3.470000 0.715000 ;
      RECT  3.270000  0.715000  3.995000 0.885000 ;
      RECT  3.270000  1.830000  3.995000 2.000000 ;
      RECT  3.270000  2.000000  3.475000 2.325000 ;
      RECT  3.640000  0.085000  3.940000 0.545000 ;
      RECT  3.645000  2.275000  3.975000 2.635000 ;
      RECT  3.735000  0.885000  3.995000 1.830000 ;
      RECT  4.110000  0.255000  4.335000 0.585000 ;
      RECT  4.145000  2.135000  4.440000 2.465000 ;
      RECT  4.165000  0.585000  4.335000 1.090000 ;
      RECT  4.165000  1.090000  4.490000 1.420000 ;
      RECT  4.165000  1.420000  4.440000 2.135000 ;
      RECT  4.505000  0.255000  4.885000 0.920000 ;
      RECT  4.665000  1.590000  4.970000 1.615000 ;
      RECT  4.665000  1.615000  4.890000 2.465000 ;
      RECT  4.715000  0.920000  4.885000 1.445000 ;
      RECT  4.715000  1.445000  4.970000 1.590000 ;
      RECT  5.055000  0.255000  5.450000 1.225000 ;
      RECT  5.055000  1.225000  7.705000 1.275000 ;
      RECT  5.060000  2.135000  5.805000 2.465000 ;
      RECT  5.140000  1.275000  6.475000 1.395000 ;
      RECT  5.205000  1.575000  5.465000 1.955000 ;
      RECT  5.620000  0.635000  6.550000 0.805000 ;
      RECT  5.620000  0.805000  6.015000 1.015000 ;
      RECT  5.635000  1.395000  5.805000 2.135000 ;
      RECT  5.665000  0.085000  6.165000 0.465000 ;
      RECT  5.975000  1.575000  6.145000 1.935000 ;
      RECT  5.975000  1.935000  6.820000 2.105000 ;
      RECT  6.000000  2.275000  6.330000 2.635000 ;
      RECT  6.305000  0.975000  7.705000 1.225000 ;
      RECT  6.335000  0.255000  6.550000 0.635000 ;
      RECT  6.605000  2.105000  6.820000 2.450000 ;
      RECT  6.720000  0.085000  7.705000 0.805000 ;
      RECT  7.060000  2.125000  8.015000 2.635000 ;
      RECT  7.355000  1.275000  7.705000 1.325000 ;
      RECT  7.385000  1.705000  8.055000 1.955000 ;
      RECT  7.885000  0.695000  9.085000 0.895000 ;
      RECT  7.885000  0.895000  8.055000 1.705000 ;
      RECT  8.185000  2.125000  8.990000 2.460000 ;
      RECT  8.420000  1.075000  8.650000 1.905000 ;
      RECT  8.465000  0.275000  9.855000 0.515000 ;
      RECT  8.820000  1.895000 10.430000 2.065000 ;
      RECT  8.820000  2.065000  8.990000 2.125000 ;
      RECT  8.830000  0.895000  9.085000 1.265000 ;
      RECT  9.160000  2.235000  9.490000 2.635000 ;
      RECT  9.285000  0.855000  9.515000 1.185000 ;
      RECT  9.285000  1.185000 10.910000 1.355000 ;
      RECT  9.660000  2.065000  9.930000 2.450000 ;
      RECT  9.685000  0.515000  9.855000 0.845000 ;
      RECT  9.685000  0.845000 10.560000 1.015000 ;
      RECT 10.035000  0.085000 10.285000 0.545000 ;
      RECT 10.100000  2.235000 10.430000 2.635000 ;
      RECT 10.105000  1.525000 10.430000 1.895000 ;
      RECT 10.465000  0.255000 10.910000 0.585000 ;
      RECT 10.600000  1.355000 10.845000 2.465000 ;
      RECT 10.730000  0.585000 10.910000 1.185000 ;
      RECT 11.080000  1.485000 11.290000 2.635000 ;
      RECT 11.120000  0.085000 11.290000 0.885000 ;
      RECT 12.025000  0.085000 12.315000 0.885000 ;
      RECT 12.025000  1.485000 12.315000 2.635000 ;
      RECT 12.530000  0.255000 12.715000 0.995000 ;
      RECT 12.530000  0.995000 13.345000 1.325000 ;
      RECT 12.530000  1.325000 12.715000 2.465000 ;
      RECT 12.885000  0.085000 13.240000 0.825000 ;
      RECT 12.885000  1.635000 13.240000 2.635000 ;
      RECT 13.910000  0.085000 14.175000 0.885000 ;
      RECT 13.910000  1.485000 14.175000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  1.445000  1.695000 1.615000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  1.785000  3.995000 1.955000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  1.105000  4.455000 1.275000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.800000  1.445000  4.970000 1.615000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.260000  1.785000  5.430000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.560000  1.785000  7.730000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.480000  1.105000  8.650000 1.275000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
    LAYER met1 ;
      RECT 1.465000 1.415000 1.755000 1.460000 ;
      RECT 1.465000 1.460000 5.030000 1.600000 ;
      RECT 1.465000 1.600000 1.755000 1.645000 ;
      RECT 3.765000 1.755000 4.055000 1.800000 ;
      RECT 3.765000 1.800000 7.790000 1.940000 ;
      RECT 3.765000 1.940000 4.055000 1.985000 ;
      RECT 4.225000 1.075000 4.515000 1.120000 ;
      RECT 4.225000 1.120000 8.710000 1.260000 ;
      RECT 4.225000 1.260000 4.515000 1.305000 ;
      RECT 4.740000 1.415000 5.030000 1.460000 ;
      RECT 4.740000 1.600000 5.030000 1.645000 ;
      RECT 5.200000 1.755000 5.490000 1.800000 ;
      RECT 5.200000 1.940000 5.490000 1.985000 ;
      RECT 7.500000 1.755000 7.790000 1.800000 ;
      RECT 7.500000 1.940000 7.790000 1.985000 ;
      RECT 8.420000 1.075000 8.710000 1.120000 ;
      RECT 8.420000 1.260000 8.710000 1.305000 ;
  END
END sky130_fd_sc_hd__sdfsbp_2
MACRO sky130_fd_sc_hd__sdfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfstp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.42000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.765000 1.335000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.995000 0.275000 12.335000 0.825000 ;
        RECT 11.995000 1.495000 12.335000 2.450000 ;
        RECT 12.145000 0.825000 12.335000 1.495000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.340000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 0.765000 0.820000 1.675000 ;
      LAYER mcon ;
        RECT 0.605000 1.105000 0.775000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.370000 1.075000 2.700000 1.600000 ;
      LAYER mcon ;
        RECT 2.445000 1.105000 2.615000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.545000 1.075000 0.835000 1.120000 ;
        RECT 0.545000 1.120000 2.675000 1.260000 ;
        RECT 0.545000 1.260000 0.835000 1.305000 ;
        RECT 2.385000 1.075000 2.675000 1.120000 ;
        RECT 2.385000 1.260000 2.675000 1.305000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 1.445000 7.065000 1.765000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.880000 1.425000 9.135000 1.545000 ;
        RECT 8.880000 1.545000 9.945000 1.725000 ;
      LAYER mcon ;
        RECT 8.940000 1.445000 9.110000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.580000 1.415000 6.870000 1.460000 ;
        RECT 6.580000 1.460000 9.170000 1.600000 ;
        RECT 6.580000 1.600000 6.870000 1.645000 ;
        RECT 8.880000 1.415000 9.170000 1.460000 ;
        RECT 8.880000 1.600000 9.170000 1.645000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.725000 3.100000 1.055000 ;
        RECT 2.905000 1.055000 3.565000 1.615000 ;
        RECT 2.905000 1.615000 3.085000 1.960000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.420000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.610000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.420000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.420000 0.085000 ;
      RECT  0.000000  2.635000 12.420000 2.805000 ;
      RECT  0.085000  0.085000  0.700000 0.595000 ;
      RECT  0.085000  1.845000  1.125000 2.025000 ;
      RECT  0.085000  2.025000  0.345000 2.465000 ;
      RECT  0.515000  2.195000  0.785000 2.635000 ;
      RECT  0.870000  0.255000  1.625000 0.555000 ;
      RECT  0.870000  0.555000  1.640000 0.575000 ;
      RECT  0.870000  0.575000  1.650000 0.595000 ;
      RECT  0.955000  2.025000  1.125000 2.255000 ;
      RECT  0.955000  2.255000  2.045000 2.465000 ;
      RECT  1.295000  1.845000  1.695000 2.085000 ;
      RECT  1.380000  0.595000  1.660000 0.600000 ;
      RECT  1.395000  0.600000  1.660000 0.605000 ;
      RECT  1.405000  0.605000  1.660000 0.610000 ;
      RECT  1.420000  0.610000  1.660000 0.615000 ;
      RECT  1.430000  0.615000  1.660000 0.620000 ;
      RECT  1.440000  0.620000  1.665000 0.630000 ;
      RECT  1.445000  0.630000  1.665000 0.635000 ;
      RECT  1.460000  0.635000  1.665000 0.645000 ;
      RECT  1.475000  0.645000  1.670000 0.660000 ;
      RECT  1.475000  0.660000  1.675000 0.665000 ;
      RECT  1.495000  0.665000  1.675000 0.705000 ;
      RECT  1.505000  0.705000  1.675000 0.710000 ;
      RECT  1.505000  0.710000  1.695000 1.845000 ;
      RECT  1.825000  0.085000  2.090000 0.545000 ;
      RECT  1.865000  0.715000  2.520000 0.905000 ;
      RECT  1.865000  0.905000  2.200000 1.770000 ;
      RECT  1.865000  1.770000  2.520000 2.085000 ;
      RECT  2.260000  0.255000  2.520000 0.715000 ;
      RECT  2.270000  2.085000  2.520000 2.465000 ;
      RECT  2.690000  0.085000  3.100000 0.555000 ;
      RECT  2.690000  2.140000  2.985000 2.635000 ;
      RECT  3.255000  1.830000  3.995000 1.990000 ;
      RECT  3.255000  1.990000  3.985000 2.000000 ;
      RECT  3.255000  2.000000  3.425000 2.325000 ;
      RECT  3.270000  0.255000  3.455000 0.715000 ;
      RECT  3.270000  0.715000  3.995000 0.885000 ;
      RECT  3.595000  2.275000  3.925000 2.635000 ;
      RECT  3.625000  0.085000  3.955000 0.545000 ;
      RECT  3.735000  0.885000  3.995000 1.830000 ;
      RECT  4.095000  2.135000  4.440000 2.465000 ;
      RECT  4.125000  0.255000  4.335000 0.585000 ;
      RECT  4.165000  0.585000  4.335000 1.090000 ;
      RECT  4.165000  1.090000  4.490000 1.420000 ;
      RECT  4.165000  1.420000  4.440000 2.135000 ;
      RECT  4.505000  0.255000  4.830000 0.920000 ;
      RECT  4.615000  1.590000  4.915000 1.615000 ;
      RECT  4.615000  1.615000  4.830000 2.465000 ;
      RECT  4.660000  0.920000  4.830000 1.445000 ;
      RECT  4.660000  1.445000  4.915000 1.590000 ;
      RECT  5.000000  0.255000  5.440000 1.225000 ;
      RECT  5.000000  1.225000  7.715000 1.275000 ;
      RECT  5.035000  2.135000  5.755000 2.465000 ;
      RECT  5.085000  1.275000  6.475000 1.395000 ;
      RECT  5.205000  1.575000  5.415000 1.955000 ;
      RECT  5.585000  1.395000  5.755000 2.135000 ;
      RECT  5.610000  0.085000  6.095000 0.465000 ;
      RECT  5.645000  0.635000  6.535000 0.805000 ;
      RECT  5.645000  0.805000  5.975000 1.015000 ;
      RECT  5.925000  1.575000  6.095000 1.935000 ;
      RECT  5.925000  1.935000  6.820000 2.105000 ;
      RECT  5.945000  2.275000  6.330000 2.635000 ;
      RECT  6.285000  0.255000  6.535000 0.635000 ;
      RECT  6.305000  0.975000  7.715000 1.225000 ;
      RECT  6.605000  2.105000  6.820000 2.450000 ;
      RECT  6.705000  0.085000  7.715000 0.805000 ;
      RECT  7.060000  2.125000  8.015000 2.635000 ;
      RECT  7.235000  1.670000  8.135000 1.955000 ;
      RECT  7.355000  1.275000  7.715000 1.325000 ;
      RECT  7.885000  0.720000  9.105000 0.905000 ;
      RECT  7.885000  0.905000  8.135000 1.670000 ;
      RECT  8.185000  2.125000  8.990000 2.460000 ;
      RECT  8.425000  1.075000  8.650000 1.905000 ;
      RECT  8.465000  0.275000  9.910000 0.545000 ;
      RECT  8.820000  0.905000  9.105000 1.255000 ;
      RECT  8.820000  1.895000 10.485000 2.065000 ;
      RECT  8.820000  2.065000  8.990000 2.125000 ;
      RECT  9.160000  2.235000  9.490000 2.635000 ;
      RECT  9.320000  0.855000  9.530000 1.195000 ;
      RECT  9.320000  1.195000 10.915000 1.365000 ;
      RECT  9.660000  2.065000  9.965000 2.450000 ;
      RECT  9.710000  0.545000  9.910000 0.785000 ;
      RECT  9.710000  0.785000 10.515000 1.015000 ;
      RECT 10.115000  0.085000 10.365000 0.545000 ;
      RECT 10.155000  1.605000 10.485000 1.895000 ;
      RECT 10.155000  2.235000 10.485000 2.635000 ;
      RECT 10.575000  0.255000 10.915000 0.585000 ;
      RECT 10.655000  1.365000 10.915000 2.465000 ;
      RECT 10.685000  0.585000 10.915000 1.195000 ;
      RECT 11.085000  0.255000 11.345000 0.995000 ;
      RECT 11.085000  0.995000 11.975000 1.325000 ;
      RECT 11.085000  1.325000 11.345000 2.465000 ;
      RECT 11.515000  0.085000 11.825000 0.825000 ;
      RECT 11.515000  1.790000 11.825000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  1.445000  1.695000 1.615000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  1.785000  3.995000 1.955000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  1.105000  4.455000 1.275000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.445000  4.915000 1.615000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.560000  1.785000  7.730000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.480000  1.105000  8.650000 1.275000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
    LAYER met1 ;
      RECT 1.465000 1.415000 1.755000 1.460000 ;
      RECT 1.465000 1.460000 4.975000 1.600000 ;
      RECT 1.465000 1.600000 1.755000 1.645000 ;
      RECT 3.765000 1.755000 4.055000 1.800000 ;
      RECT 3.765000 1.800000 7.790000 1.940000 ;
      RECT 3.765000 1.940000 4.055000 1.985000 ;
      RECT 4.225000 1.075000 4.515000 1.120000 ;
      RECT 4.225000 1.120000 8.710000 1.260000 ;
      RECT 4.225000 1.260000 4.515000 1.305000 ;
      RECT 4.685000 1.415000 4.975000 1.460000 ;
      RECT 4.685000 1.600000 4.975000 1.645000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 7.500000 1.755000 7.790000 1.800000 ;
      RECT 7.500000 1.940000 7.790000 1.985000 ;
      RECT 8.420000 1.075000 8.710000 1.120000 ;
      RECT 8.420000 1.260000 8.710000 1.305000 ;
  END
END sky130_fd_sc_hd__sdfstp_1
MACRO sky130_fd_sc_hd__sdfstp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfstp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.88000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.765000 1.335000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.519750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.035000 0.255000 12.365000 0.825000 ;
        RECT 12.035000 1.495000 12.365000 2.450000 ;
        RECT 12.145000 0.825000 12.365000 1.495000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.340000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 0.765000 0.820000 1.675000 ;
      LAYER mcon ;
        RECT 0.605000 1.105000 0.775000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.370000 1.075000 2.700000 1.600000 ;
      LAYER mcon ;
        RECT 2.445000 1.105000 2.615000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.545000 1.075000 0.835000 1.120000 ;
        RECT 0.545000 1.120000 2.675000 1.260000 ;
        RECT 0.545000 1.260000 0.835000 1.305000 ;
        RECT 2.385000 1.075000 2.675000 1.120000 ;
        RECT 2.385000 1.260000 2.675000 1.305000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 1.445000 7.065000 1.765000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.880000 1.425000 9.135000 1.545000 ;
        RECT 8.880000 1.545000 9.945000 1.725000 ;
      LAYER mcon ;
        RECT 8.940000 1.445000 9.110000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.580000 1.415000 6.870000 1.460000 ;
        RECT 6.580000 1.460000 9.170000 1.600000 ;
        RECT 6.580000 1.600000 6.870000 1.645000 ;
        RECT 8.880000 1.415000 9.170000 1.460000 ;
        RECT 8.880000 1.600000 9.170000 1.645000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.725000 3.100000 1.055000 ;
        RECT 2.905000 1.055000 3.565000 1.615000 ;
        RECT 2.905000 1.615000 3.085000 1.960000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.880000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 13.070000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.880000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.880000 0.085000 ;
      RECT  0.000000  2.635000 12.880000 2.805000 ;
      RECT  0.085000  0.085000  0.700000 0.595000 ;
      RECT  0.085000  1.845000  1.125000 2.025000 ;
      RECT  0.085000  2.025000  0.345000 2.465000 ;
      RECT  0.515000  2.195000  0.785000 2.635000 ;
      RECT  0.870000  0.255000  1.625000 0.555000 ;
      RECT  0.870000  0.555000  1.640000 0.575000 ;
      RECT  0.870000  0.575000  1.650000 0.595000 ;
      RECT  0.955000  2.025000  1.125000 2.255000 ;
      RECT  0.955000  2.255000  2.045000 2.465000 ;
      RECT  1.295000  1.845000  1.695000 2.085000 ;
      RECT  1.380000  0.595000  1.660000 0.600000 ;
      RECT  1.395000  0.600000  1.660000 0.605000 ;
      RECT  1.405000  0.605000  1.660000 0.610000 ;
      RECT  1.420000  0.610000  1.660000 0.615000 ;
      RECT  1.430000  0.615000  1.660000 0.620000 ;
      RECT  1.440000  0.620000  1.665000 0.630000 ;
      RECT  1.445000  0.630000  1.665000 0.635000 ;
      RECT  1.460000  0.635000  1.665000 0.645000 ;
      RECT  1.475000  0.645000  1.670000 0.660000 ;
      RECT  1.475000  0.660000  1.675000 0.665000 ;
      RECT  1.495000  0.665000  1.675000 0.705000 ;
      RECT  1.505000  0.705000  1.675000 0.710000 ;
      RECT  1.505000  0.710000  1.695000 1.845000 ;
      RECT  1.825000  0.085000  2.090000 0.545000 ;
      RECT  1.865000  0.715000  2.520000 0.905000 ;
      RECT  1.865000  0.905000  2.200000 1.770000 ;
      RECT  1.865000  1.770000  2.520000 2.085000 ;
      RECT  2.260000  0.255000  2.520000 0.715000 ;
      RECT  2.270000  2.085000  2.520000 2.465000 ;
      RECT  2.690000  0.085000  3.100000 0.555000 ;
      RECT  2.690000  2.140000  2.985000 2.635000 ;
      RECT  3.255000  1.830000  3.995000 1.990000 ;
      RECT  3.255000  1.990000  3.985000 2.000000 ;
      RECT  3.255000  2.000000  3.425000 2.325000 ;
      RECT  3.270000  0.255000  3.455000 0.715000 ;
      RECT  3.270000  0.715000  3.995000 0.885000 ;
      RECT  3.595000  2.275000  3.925000 2.635000 ;
      RECT  3.625000  0.085000  3.955000 0.545000 ;
      RECT  3.735000  0.885000  3.995000 1.830000 ;
      RECT  4.095000  2.135000  4.440000 2.465000 ;
      RECT  4.125000  0.255000  4.335000 0.585000 ;
      RECT  4.165000  0.585000  4.335000 1.090000 ;
      RECT  4.165000  1.090000  4.490000 1.420000 ;
      RECT  4.165000  1.420000  4.440000 2.135000 ;
      RECT  4.505000  0.255000  4.830000 0.920000 ;
      RECT  4.615000  1.590000  4.915000 1.615000 ;
      RECT  4.615000  1.615000  4.830000 2.465000 ;
      RECT  4.660000  0.920000  4.830000 1.445000 ;
      RECT  4.660000  1.445000  4.915000 1.590000 ;
      RECT  5.000000  0.255000  5.440000 1.225000 ;
      RECT  5.000000  1.225000  7.715000 1.275000 ;
      RECT  5.035000  2.135000  5.755000 2.465000 ;
      RECT  5.085000  1.275000  6.475000 1.395000 ;
      RECT  5.205000  1.575000  5.415000 1.955000 ;
      RECT  5.585000  1.395000  5.755000 2.135000 ;
      RECT  5.610000  0.085000  6.095000 0.465000 ;
      RECT  5.645000  0.635000  6.535000 0.805000 ;
      RECT  5.645000  0.805000  5.975000 1.015000 ;
      RECT  5.925000  1.575000  6.095000 1.935000 ;
      RECT  5.925000  1.935000  6.820000 2.105000 ;
      RECT  5.945000  2.275000  6.330000 2.635000 ;
      RECT  6.285000  0.255000  6.535000 0.635000 ;
      RECT  6.305000  0.975000  7.715000 1.225000 ;
      RECT  6.605000  2.105000  6.820000 2.450000 ;
      RECT  6.705000  0.085000  7.715000 0.805000 ;
      RECT  7.060000  2.125000  8.015000 2.635000 ;
      RECT  7.235000  1.670000  8.135000 1.955000 ;
      RECT  7.355000  1.275000  7.715000 1.325000 ;
      RECT  7.885000  0.720000  9.105000 0.905000 ;
      RECT  7.885000  0.905000  8.135000 1.670000 ;
      RECT  8.185000  2.125000  8.990000 2.460000 ;
      RECT  8.425000  1.075000  8.650000 1.905000 ;
      RECT  8.465000  0.275000  9.910000 0.545000 ;
      RECT  8.820000  0.905000  9.105000 1.255000 ;
      RECT  8.820000  1.895000 10.485000 2.065000 ;
      RECT  8.820000  2.065000  8.990000 2.125000 ;
      RECT  9.160000  2.235000  9.490000 2.635000 ;
      RECT  9.320000  0.855000  9.530000 1.195000 ;
      RECT  9.320000  1.195000 10.915000 1.365000 ;
      RECT  9.660000  2.065000  9.965000 2.450000 ;
      RECT  9.710000  0.545000  9.910000 0.785000 ;
      RECT  9.710000  0.785000 10.515000 1.015000 ;
      RECT 10.115000  0.085000 10.365000 0.545000 ;
      RECT 10.155000  1.605000 10.485000 1.895000 ;
      RECT 10.155000  2.235000 10.485000 2.635000 ;
      RECT 10.575000  0.255000 10.915000 0.585000 ;
      RECT 10.655000  1.365000 10.915000 2.465000 ;
      RECT 10.685000  0.585000 10.915000 1.195000 ;
      RECT 11.085000  0.255000 11.345000 0.995000 ;
      RECT 11.085000  0.995000 11.975000 1.325000 ;
      RECT 11.085000  1.325000 11.345000 2.465000 ;
      RECT 11.570000  0.085000 11.865000 0.825000 ;
      RECT 11.570000  1.790000 11.820000 2.635000 ;
      RECT 12.535000  0.085000 12.795000 0.885000 ;
      RECT 12.535000  1.495000 12.795000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  1.445000  1.695000 1.615000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  1.785000  3.995000 1.955000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  1.105000  4.455000 1.275000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.445000  4.915000 1.615000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.560000  1.785000  7.730000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.480000  1.105000  8.650000 1.275000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
    LAYER met1 ;
      RECT 1.465000 1.415000 1.755000 1.460000 ;
      RECT 1.465000 1.460000 4.975000 1.600000 ;
      RECT 1.465000 1.600000 1.755000 1.645000 ;
      RECT 3.765000 1.755000 4.055000 1.800000 ;
      RECT 3.765000 1.800000 7.790000 1.940000 ;
      RECT 3.765000 1.940000 4.055000 1.985000 ;
      RECT 4.225000 1.075000 4.515000 1.120000 ;
      RECT 4.225000 1.120000 8.710000 1.260000 ;
      RECT 4.225000 1.260000 4.515000 1.305000 ;
      RECT 4.685000 1.415000 4.975000 1.460000 ;
      RECT 4.685000 1.600000 4.975000 1.645000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 7.500000 1.755000 7.790000 1.800000 ;
      RECT 7.500000 1.940000 7.790000 1.985000 ;
      RECT 8.420000 1.075000 8.710000 1.120000 ;
      RECT 8.420000 1.260000 8.710000 1.305000 ;
  END
END sky130_fd_sc_hd__sdfstp_2
MACRO sky130_fd_sc_hd__sdfstp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfstp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.80000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.765000 1.335000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.040000 0.275000 12.370000 0.825000 ;
        RECT 12.040000 1.495000 12.370000 2.450000 ;
        RECT 12.145000 0.825000 12.370000 1.055000 ;
        RECT 12.145000 1.055000 13.210000 1.325000 ;
        RECT 12.145000 1.325000 12.370000 1.495000 ;
        RECT 12.880000 0.255000 13.210000 1.055000 ;
        RECT 12.880000 1.325000 13.210000 2.465000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.340000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 0.765000 0.820000 1.675000 ;
      LAYER mcon ;
        RECT 0.605000 1.105000 0.775000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.370000 1.075000 2.700000 1.600000 ;
      LAYER mcon ;
        RECT 2.445000 1.105000 2.615000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.545000 1.075000 0.835000 1.120000 ;
        RECT 0.545000 1.120000 2.675000 1.260000 ;
        RECT 0.545000 1.260000 0.835000 1.305000 ;
        RECT 2.385000 1.075000 2.675000 1.120000 ;
        RECT 2.385000 1.260000 2.675000 1.305000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 1.445000 7.065000 1.765000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.880000 1.425000 9.135000 1.545000 ;
        RECT 8.880000 1.545000 9.945000 1.725000 ;
      LAYER mcon ;
        RECT 8.940000 1.445000 9.110000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.580000 1.415000 6.870000 1.460000 ;
        RECT 6.580000 1.460000 9.170000 1.600000 ;
        RECT 6.580000 1.600000 6.870000 1.645000 ;
        RECT 8.880000 1.415000 9.170000 1.460000 ;
        RECT 8.880000 1.600000 9.170000 1.645000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.725000 3.100000 1.055000 ;
        RECT 2.905000 1.055000 3.565000 1.615000 ;
        RECT 2.905000 1.615000 3.085000 1.960000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.800000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 13.990000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.800000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.800000 0.085000 ;
      RECT  0.000000  2.635000 13.800000 2.805000 ;
      RECT  0.085000  0.085000  0.700000 0.595000 ;
      RECT  0.085000  1.845000  1.125000 2.025000 ;
      RECT  0.085000  2.025000  0.345000 2.465000 ;
      RECT  0.515000  2.195000  0.785000 2.635000 ;
      RECT  0.870000  0.255000  1.625000 0.555000 ;
      RECT  0.870000  0.555000  1.640000 0.575000 ;
      RECT  0.870000  0.575000  1.650000 0.595000 ;
      RECT  0.955000  2.025000  1.125000 2.255000 ;
      RECT  0.955000  2.255000  2.045000 2.465000 ;
      RECT  1.295000  1.845000  1.695000 2.085000 ;
      RECT  1.380000  0.595000  1.660000 0.600000 ;
      RECT  1.395000  0.600000  1.660000 0.605000 ;
      RECT  1.405000  0.605000  1.660000 0.610000 ;
      RECT  1.420000  0.610000  1.660000 0.615000 ;
      RECT  1.430000  0.615000  1.660000 0.620000 ;
      RECT  1.440000  0.620000  1.665000 0.630000 ;
      RECT  1.445000  0.630000  1.665000 0.635000 ;
      RECT  1.460000  0.635000  1.665000 0.645000 ;
      RECT  1.475000  0.645000  1.670000 0.660000 ;
      RECT  1.475000  0.660000  1.675000 0.665000 ;
      RECT  1.495000  0.665000  1.675000 0.705000 ;
      RECT  1.505000  0.705000  1.675000 0.710000 ;
      RECT  1.505000  0.710000  1.695000 1.845000 ;
      RECT  1.825000  0.085000  2.090000 0.545000 ;
      RECT  1.865000  0.715000  2.520000 0.905000 ;
      RECT  1.865000  0.905000  2.200000 1.770000 ;
      RECT  1.865000  1.770000  2.520000 2.085000 ;
      RECT  2.260000  0.255000  2.520000 0.715000 ;
      RECT  2.270000  2.085000  2.520000 2.465000 ;
      RECT  2.690000  0.085000  3.100000 0.555000 ;
      RECT  2.690000  2.140000  2.985000 2.635000 ;
      RECT  3.255000  1.830000  3.995000 1.990000 ;
      RECT  3.255000  1.990000  3.985000 2.000000 ;
      RECT  3.255000  2.000000  3.425000 2.325000 ;
      RECT  3.270000  0.255000  3.455000 0.715000 ;
      RECT  3.270000  0.715000  3.995000 0.885000 ;
      RECT  3.595000  2.275000  3.925000 2.635000 ;
      RECT  3.625000  0.085000  3.955000 0.545000 ;
      RECT  3.735000  0.885000  3.995000 1.830000 ;
      RECT  4.095000  2.135000  4.440000 2.465000 ;
      RECT  4.125000  0.255000  4.335000 0.585000 ;
      RECT  4.165000  0.585000  4.335000 1.090000 ;
      RECT  4.165000  1.090000  4.490000 1.420000 ;
      RECT  4.165000  1.420000  4.440000 2.135000 ;
      RECT  4.505000  0.255000  4.830000 0.920000 ;
      RECT  4.615000  1.590000  4.915000 1.615000 ;
      RECT  4.615000  1.615000  4.830000 2.465000 ;
      RECT  4.660000  0.920000  4.830000 1.445000 ;
      RECT  4.660000  1.445000  4.915000 1.590000 ;
      RECT  5.000000  0.255000  5.440000 1.225000 ;
      RECT  5.000000  1.225000  7.715000 1.275000 ;
      RECT  5.035000  2.135000  5.755000 2.465000 ;
      RECT  5.085000  1.275000  6.475000 1.395000 ;
      RECT  5.205000  1.575000  5.415000 1.955000 ;
      RECT  5.585000  1.395000  5.755000 2.135000 ;
      RECT  5.610000  0.085000  6.095000 0.465000 ;
      RECT  5.645000  0.635000  6.535000 0.805000 ;
      RECT  5.645000  0.805000  5.975000 1.015000 ;
      RECT  5.925000  1.575000  6.095000 1.935000 ;
      RECT  5.925000  1.935000  6.820000 2.105000 ;
      RECT  5.945000  2.275000  6.330000 2.635000 ;
      RECT  6.285000  0.255000  6.535000 0.635000 ;
      RECT  6.305000  0.975000  7.715000 1.225000 ;
      RECT  6.605000  2.105000  6.820000 2.450000 ;
      RECT  6.705000  0.085000  7.715000 0.805000 ;
      RECT  7.060000  2.125000  8.015000 2.635000 ;
      RECT  7.235000  1.670000  8.135000 1.955000 ;
      RECT  7.355000  1.275000  7.715000 1.325000 ;
      RECT  7.885000  0.720000  9.105000 0.905000 ;
      RECT  7.885000  0.905000  8.135000 1.670000 ;
      RECT  8.185000  2.125000  8.990000 2.460000 ;
      RECT  8.425000  1.075000  8.650000 1.905000 ;
      RECT  8.465000  0.275000  9.910000 0.545000 ;
      RECT  8.820000  0.905000  9.105000 1.255000 ;
      RECT  8.820000  1.895000 10.485000 2.065000 ;
      RECT  8.820000  2.065000  8.990000 2.125000 ;
      RECT  9.160000  2.235000  9.490000 2.635000 ;
      RECT  9.320000  0.855000  9.530000 1.195000 ;
      RECT  9.320000  1.195000 10.915000 1.365000 ;
      RECT  9.660000  2.065000  9.965000 2.450000 ;
      RECT  9.710000  0.545000  9.910000 0.785000 ;
      RECT  9.710000  0.785000 10.515000 1.015000 ;
      RECT 10.115000  0.085000 10.365000 0.545000 ;
      RECT 10.155000  1.605000 10.485000 1.895000 ;
      RECT 10.155000  2.235000 10.485000 2.635000 ;
      RECT 10.575000  0.255000 10.915000 0.585000 ;
      RECT 10.655000  1.365000 10.915000 2.465000 ;
      RECT 10.685000  0.585000 10.915000 1.195000 ;
      RECT 11.085000  0.255000 11.345000 0.995000 ;
      RECT 11.085000  0.995000 11.975000 1.325000 ;
      RECT 11.085000  1.325000 11.345000 2.465000 ;
      RECT 11.515000  0.085000 11.870000 0.825000 ;
      RECT 11.515000  1.495000 11.870000 2.635000 ;
      RECT 12.540000  0.085000 12.710000 0.885000 ;
      RECT 12.540000  1.495000 12.710000 2.635000 ;
      RECT 13.380000  0.085000 13.715000 0.885000 ;
      RECT 13.380000  1.495000 13.715000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  1.445000  1.695000 1.615000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  1.785000  3.995000 1.955000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  1.105000  4.455000 1.275000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.445000  4.915000 1.615000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.560000  1.785000  7.730000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.480000  1.105000  8.650000 1.275000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
    LAYER met1 ;
      RECT 1.465000 1.415000 1.755000 1.460000 ;
      RECT 1.465000 1.460000 4.975000 1.600000 ;
      RECT 1.465000 1.600000 1.755000 1.645000 ;
      RECT 3.765000 1.755000 4.055000 1.800000 ;
      RECT 3.765000 1.800000 7.790000 1.940000 ;
      RECT 3.765000 1.940000 4.055000 1.985000 ;
      RECT 4.225000 1.075000 4.515000 1.120000 ;
      RECT 4.225000 1.120000 8.710000 1.260000 ;
      RECT 4.225000 1.260000 4.515000 1.305000 ;
      RECT 4.685000 1.415000 4.975000 1.460000 ;
      RECT 4.685000 1.600000 4.975000 1.645000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 7.500000 1.755000 7.790000 1.800000 ;
      RECT 7.500000 1.940000 7.790000 1.985000 ;
      RECT 8.420000 1.075000 8.710000 1.120000 ;
      RECT 8.420000 1.260000 8.710000 1.305000 ;
  END
END sky130_fd_sc_hd__sdfstp_4
MACRO sky130_fd_sc_hd__sdfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.440000 1.355000 2.775000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.180000 0.305000 9.530000 0.725000 ;
        RECT 9.180000 0.725000 9.560000 0.790000 ;
        RECT 9.180000 0.790000 9.610000 0.825000 ;
        RECT 9.200000 1.505000 9.610000 1.540000 ;
        RECT 9.200000 1.540000 9.530000 2.465000 ;
        RECT 9.355000 1.430000 9.610000 1.505000 ;
        RECT 9.390000 0.825000 9.610000 1.430000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.685000 0.265000 10.940000 0.795000 ;
        RECT 10.685000 1.445000 10.940000 2.325000 ;
        RECT 10.730000 0.795000 10.940000 1.445000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.515000 1.055000 3.995000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.760000 0.750000 3.235000 0.785000 ;
        RECT 1.760000 0.785000 2.010000 0.810000 ;
        RECT 1.760000 0.810000 1.990000 0.820000 ;
        RECT 1.760000 0.820000 1.975000 0.835000 ;
        RECT 1.760000 0.835000 1.970000 0.840000 ;
        RECT 1.760000 0.840000 1.965000 0.850000 ;
        RECT 1.760000 0.850000 1.960000 0.855000 ;
        RECT 1.760000 0.855000 1.955000 0.860000 ;
        RECT 1.760000 0.860000 1.950000 0.870000 ;
        RECT 1.760000 0.870000 1.945000 0.875000 ;
        RECT 1.760000 0.875000 1.940000 0.880000 ;
        RECT 1.760000 0.880000 1.930000 1.685000 ;
        RECT 1.790000 0.735000 3.235000 0.750000 ;
        RECT 1.805000 0.725000 3.235000 0.735000 ;
        RECT 1.820000 0.715000 3.235000 0.725000 ;
        RECT 1.830000 0.705000 3.235000 0.715000 ;
        RECT 1.840000 0.690000 3.235000 0.705000 ;
        RECT 1.860000 0.655000 3.235000 0.690000 ;
        RECT 1.875000 0.615000 3.235000 0.655000 ;
        RECT 2.455000 0.305000 2.630000 0.615000 ;
        RECT 3.065000 0.785000 3.235000 1.115000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.810000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.810000 0.970000 ;
      RECT  0.615000  0.970000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.420000  0.255000  1.705000 0.585000 ;
      RECT  1.420000  0.585000  1.590000 1.860000 ;
      RECT  1.420000  1.860000  3.230000 2.075000 ;
      RECT  1.420000  2.075000  1.705000 2.445000 ;
      RECT  1.875000  2.245000  2.205000 2.635000 ;
      RECT  1.955000  0.085000  2.285000 0.445000 ;
      RECT  2.100000  0.955000  2.445000 1.125000 ;
      RECT  2.100000  1.125000  2.270000 1.860000 ;
      RECT  2.675000  2.245000  3.570000 2.415000 ;
      RECT  2.800000  0.275000  3.575000 0.445000 ;
      RECT  3.060000  1.355000  3.255000 1.685000 ;
      RECT  3.060000  1.685000  3.230000 1.860000 ;
      RECT  3.400000  1.825000  4.335000 1.995000 ;
      RECT  3.400000  1.995000  3.570000 2.245000 ;
      RECT  3.405000  0.445000  3.575000 0.715000 ;
      RECT  3.405000  0.715000  4.335000 0.885000 ;
      RECT  3.740000  2.165000  3.910000 2.635000 ;
      RECT  3.745000  0.085000  3.945000 0.545000 ;
      RECT  4.165000  0.365000  4.515000 0.535000 ;
      RECT  4.165000  0.535000  4.335000 0.715000 ;
      RECT  4.165000  0.885000  4.335000 1.825000 ;
      RECT  4.165000  1.995000  4.335000 2.070000 ;
      RECT  4.165000  2.070000  4.450000 2.440000 ;
      RECT  4.505000  0.705000  5.085000 1.035000 ;
      RECT  4.505000  1.035000  4.745000 1.905000 ;
      RECT  4.645000  2.190000  5.715000 2.360000 ;
      RECT  4.685000  0.365000  5.425000 0.535000 ;
      RECT  4.935000  1.655000  5.375000 2.010000 ;
      RECT  5.255000  0.535000  5.425000 1.315000 ;
      RECT  5.255000  1.315000  6.055000 1.485000 ;
      RECT  5.545000  1.485000  6.055000 1.575000 ;
      RECT  5.545000  1.575000  5.715000 2.190000 ;
      RECT  5.595000  0.765000  6.395000 1.065000 ;
      RECT  5.595000  1.065000  5.765000 1.095000 ;
      RECT  5.675000  0.085000  6.045000 0.585000 ;
      RECT  5.885000  1.245000  6.055000 1.315000 ;
      RECT  5.885000  1.835000  6.055000 2.635000 ;
      RECT  6.225000  0.365000  6.685000 0.535000 ;
      RECT  6.225000  0.535000  6.395000 0.765000 ;
      RECT  6.225000  1.065000  6.395000 2.135000 ;
      RECT  6.225000  2.135000  6.475000 2.465000 ;
      RECT  6.565000  0.705000  7.115000 1.035000 ;
      RECT  6.565000  1.245000  6.755000 1.965000 ;
      RECT  6.700000  2.165000  7.585000 2.335000 ;
      RECT  6.915000  0.365000  7.455000 0.535000 ;
      RECT  6.925000  1.035000  7.115000 1.575000 ;
      RECT  6.925000  1.575000  7.245000 1.905000 ;
      RECT  7.285000  0.535000  7.455000 0.995000 ;
      RECT  7.285000  0.995000  8.315000 1.325000 ;
      RECT  7.285000  1.325000  7.585000 1.405000 ;
      RECT  7.415000  1.405000  7.585000 2.165000 ;
      RECT  7.700000  0.085000  8.070000 0.615000 ;
      RECT  7.755000  1.575000  8.670000 1.905000 ;
      RECT  7.765000  2.135000  8.070000 2.635000 ;
      RECT  8.340000  0.300000  8.670000 0.825000 ;
      RECT  8.380000  1.905000  8.670000 2.455000 ;
      RECT  8.485000  0.825000  8.670000 0.995000 ;
      RECT  8.485000  0.995000  9.220000 1.325000 ;
      RECT  8.485000  1.325000  8.670000 1.575000 ;
      RECT  8.840000  0.085000  9.010000 0.695000 ;
      RECT  8.840000  1.625000  9.010000 2.635000 ;
      RECT  9.700000  0.345000  9.950000 0.620000 ;
      RECT  9.700000  1.685000 10.030000 2.425000 ;
      RECT  9.780000  0.620000  9.950000 0.995000 ;
      RECT  9.780000  0.995000 10.560000 1.325000 ;
      RECT  9.780000  1.325000 10.030000 1.685000 ;
      RECT 10.185000  0.085000 10.515000 0.805000 ;
      RECT 10.210000  1.495000 10.515000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.645000  1.785000  0.815000 1.955000 ;
      RECT  1.015000  0.765000  1.185000 0.935000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  0.765000  4.915000 0.935000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.165000  1.785000  5.335000 1.955000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.575000  1.785000  6.745000 1.955000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  0.765000  6.755000 0.935000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 0.585000 1.755000 0.875000 1.800000 ;
      RECT 0.585000 1.800000 6.805000 1.940000 ;
      RECT 0.585000 1.940000 0.875000 1.985000 ;
      RECT 0.955000 0.735000 1.245000 0.780000 ;
      RECT 0.955000 0.780000 6.815000 0.920000 ;
      RECT 0.955000 0.920000 1.245000 0.965000 ;
      RECT 4.685000 0.735000 4.975000 0.780000 ;
      RECT 4.685000 0.920000 4.975000 0.965000 ;
      RECT 5.105000 1.755000 5.395000 1.800000 ;
      RECT 5.105000 1.940000 5.395000 1.985000 ;
      RECT 6.515000 1.755000 6.805000 1.800000 ;
      RECT 6.515000 1.940000 6.805000 1.985000 ;
      RECT 6.525000 0.735000 6.815000 0.780000 ;
      RECT 6.525000 0.920000 6.815000 0.965000 ;
  END
END sky130_fd_sc_hd__sdfxbp_1
MACRO sky130_fd_sc_hd__sdfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.460000 1.355000 2.795000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.255000 0.255000 9.585000 0.790000 ;
        RECT 9.255000 0.790000 9.615000 0.825000 ;
        RECT 9.255000 1.495000 9.615000 1.530000 ;
        RECT 9.255000 1.530000 9.585000 2.430000 ;
        RECT 9.410000 0.825000 9.615000 0.890000 ;
        RECT 9.410000 1.430000 9.615000 1.495000 ;
        RECT 9.445000 0.890000 9.615000 1.430000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.190000 0.265000 11.440000 0.795000 ;
        RECT 11.190000 1.445000 11.440000 2.325000 ;
        RECT 11.235000 0.795000 11.440000 1.445000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.535000 1.035000 4.035000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.780000 0.615000 3.255000 0.785000 ;
        RECT 1.780000 0.785000 1.950000 1.685000 ;
        RECT 2.475000 0.305000 2.650000 0.615000 ;
        RECT 3.085000 0.785000 3.255000 1.115000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.150000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.810000 0.805000 ;
      RECT  0.180000  1.795000  0.845000 1.965000 ;
      RECT  0.180000  1.965000  0.350000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.520000  2.135000  0.850000 2.635000 ;
      RECT  0.615000  0.805000  0.810000 0.970000 ;
      RECT  0.615000  0.970000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.245000 0.715000 ;
      RECT  1.020000  0.715000  1.245000 2.465000 ;
      RECT  1.435000  0.275000  1.805000 0.445000 ;
      RECT  1.435000  0.445000  1.605000 1.860000 ;
      RECT  1.435000  1.860000  3.250000 2.075000 ;
      RECT  1.435000  2.075000  1.710000 2.445000 ;
      RECT  1.880000  2.245000  2.210000 2.635000 ;
      RECT  1.975000  0.085000  2.305000 0.445000 ;
      RECT  2.120000  0.955000  2.465000 1.125000 ;
      RECT  2.120000  1.125000  2.290000 1.860000 ;
      RECT  2.695000  2.245000  3.590000 2.415000 ;
      RECT  2.820000  0.275000  3.595000 0.445000 ;
      RECT  3.080000  1.355000  3.275000 1.685000 ;
      RECT  3.080000  1.685000  3.250000 1.860000 ;
      RECT  3.420000  1.825000  4.375000 1.995000 ;
      RECT  3.420000  1.995000  3.590000 2.245000 ;
      RECT  3.425000  0.445000  3.595000 0.695000 ;
      RECT  3.425000  0.695000  4.375000 0.865000 ;
      RECT  3.760000  2.165000  3.930000 2.635000 ;
      RECT  3.765000  0.085000  3.965000 0.525000 ;
      RECT  4.205000  0.365000  4.555000 0.535000 ;
      RECT  4.205000  0.535000  4.375000 0.695000 ;
      RECT  4.205000  0.865000  4.375000 1.825000 ;
      RECT  4.205000  1.995000  4.375000 2.065000 ;
      RECT  4.205000  2.065000  4.485000 2.440000 ;
      RECT  4.545000  0.705000  5.125000 1.035000 ;
      RECT  4.545000  1.035000  4.785000 1.905000 ;
      RECT  4.685000  2.190000  5.755000 2.360000 ;
      RECT  4.725000  0.365000  5.465000 0.535000 ;
      RECT  4.975000  1.655000  5.415000 2.010000 ;
      RECT  5.295000  0.535000  5.465000 1.315000 ;
      RECT  5.295000  1.315000  6.095000 1.485000 ;
      RECT  5.585000  1.485000  6.095000 1.575000 ;
      RECT  5.585000  1.575000  5.755000 2.190000 ;
      RECT  5.635000  0.765000  6.435000 1.065000 ;
      RECT  5.635000  1.065000  5.805000 1.095000 ;
      RECT  5.715000  0.085000  6.085000 0.585000 ;
      RECT  5.925000  1.245000  6.095000 1.315000 ;
      RECT  5.925000  1.835000  6.095000 2.635000 ;
      RECT  6.265000  0.365000  6.725000 0.535000 ;
      RECT  6.265000  0.535000  6.435000 0.765000 ;
      RECT  6.265000  1.065000  6.435000 2.135000 ;
      RECT  6.265000  2.135000  6.515000 2.465000 ;
      RECT  6.605000  0.705000  7.155000 1.035000 ;
      RECT  6.605000  1.245000  6.795000 1.965000 ;
      RECT  6.740000  2.165000  7.625000 2.335000 ;
      RECT  6.955000  0.365000  7.495000 0.535000 ;
      RECT  6.965000  1.035000  7.155000 1.575000 ;
      RECT  6.965000  1.575000  7.285000 1.905000 ;
      RECT  7.325000  0.535000  7.495000 0.995000 ;
      RECT  7.325000  0.995000  8.370000 1.325000 ;
      RECT  7.325000  1.325000  7.625000 1.405000 ;
      RECT  7.455000  1.405000  7.625000 2.165000 ;
      RECT  7.740000  0.085000  8.110000 0.615000 ;
      RECT  7.795000  1.575000  8.725000 1.905000 ;
      RECT  7.805000  2.135000  8.110000 2.635000 ;
      RECT  8.360000  0.300000  8.725000 0.825000 ;
      RECT  8.395000  1.905000  8.725000 2.455000 ;
      RECT  8.540000  0.825000  8.725000 0.995000 ;
      RECT  8.540000  0.995000  9.275000 1.325000 ;
      RECT  8.540000  1.325000  8.725000 1.575000 ;
      RECT  8.895000  0.085000  9.085000 0.695000 ;
      RECT  8.895000  1.625000  9.075000 2.635000 ;
      RECT  9.755000  0.085000  9.985000 0.690000 ;
      RECT  9.765000  1.615000  9.935000 2.635000 ;
      RECT 10.205000  0.345000 10.455000 0.995000 ;
      RECT 10.205000  0.995000 11.065000 1.325000 ;
      RECT 10.205000  1.325000 10.535000 2.425000 ;
      RECT 10.690000  0.085000 11.020000 0.805000 ;
      RECT 10.715000  1.495000 11.020000 2.635000 ;
      RECT 11.610000  0.085000 11.780000 0.955000 ;
      RECT 11.610000  1.395000 11.780000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.645000  1.785000  0.815000 1.955000 ;
      RECT  1.050000  0.765000  1.220000 0.935000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  0.765000  4.915000 0.935000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.625000  1.785000  6.795000 1.955000 ;
      RECT  6.640000  0.765000  6.810000 0.935000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
    LAYER met1 ;
      RECT 0.585000 1.755000 0.875000 1.800000 ;
      RECT 0.585000 1.800000 6.855000 1.940000 ;
      RECT 0.585000 1.940000 0.875000 1.985000 ;
      RECT 0.990000 0.735000 1.280000 0.780000 ;
      RECT 0.990000 0.780000 6.870000 0.920000 ;
      RECT 0.990000 0.920000 1.280000 0.965000 ;
      RECT 4.685000 0.735000 4.975000 0.780000 ;
      RECT 4.685000 0.920000 4.975000 0.965000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 6.565000 1.755000 6.855000 1.800000 ;
      RECT 6.565000 1.940000 6.855000 1.985000 ;
      RECT 6.580000 0.735000 6.870000 0.780000 ;
      RECT 6.580000 0.920000 6.870000 0.965000 ;
  END
END sky130_fd_sc_hd__sdfxbp_2
MACRO sky130_fd_sc_hd__sdfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.460000 1.355000 2.790000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.230000 0.305000 9.575000 0.820000 ;
        RECT 9.230000 1.505000 9.575000 2.395000 ;
        RECT 9.405000 0.820000 9.575000 1.505000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.530000 1.055000 3.990000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.760000 0.635000 3.250000 0.785000 ;
        RECT 1.760000 0.785000 1.990000 0.835000 ;
        RECT 1.760000 0.835000 1.930000 1.685000 ;
        RECT 1.870000 0.615000 3.250000 0.635000 ;
        RECT 2.475000 0.305000 2.650000 0.615000 ;
        RECT 3.065000 0.785000 3.250000 1.095000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.810000 0.805000 ;
      RECT 0.180000  1.795000 0.845000 1.965000 ;
      RECT 0.180000  1.965000 0.350000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.520000  2.135000 0.850000 2.635000 ;
      RECT 0.615000  0.805000 0.810000 0.970000 ;
      RECT 0.615000  0.970000 0.845000 1.795000 ;
      RECT 1.015000  0.345000 1.230000 0.715000 ;
      RECT 1.020000  0.715000 1.230000 2.465000 ;
      RECT 1.420000  0.260000 1.790000 0.465000 ;
      RECT 1.420000  0.465000 1.590000 1.860000 ;
      RECT 1.420000  1.860000 3.220000 2.075000 ;
      RECT 1.420000  2.075000 1.710000 2.445000 ;
      RECT 1.880000  2.245000 2.210000 2.635000 ;
      RECT 1.960000  0.085000 2.305000 0.445000 ;
      RECT 2.115000  0.960000 2.460000 1.130000 ;
      RECT 2.115000  1.130000 2.290000 1.860000 ;
      RECT 2.690000  2.245000 3.560000 2.415000 ;
      RECT 2.820000  0.275000 3.590000 0.445000 ;
      RECT 3.050000  1.305000 3.270000 1.635000 ;
      RECT 3.050000  1.635000 3.220000 1.860000 ;
      RECT 3.390000  1.825000 4.350000 1.995000 ;
      RECT 3.390000  1.995000 3.560000 2.245000 ;
      RECT 3.420000  0.445000 3.590000 0.715000 ;
      RECT 3.420000  0.715000 4.350000 0.885000 ;
      RECT 3.730000  2.165000 3.925000 2.635000 ;
      RECT 3.760000  0.085000 3.960000 0.545000 ;
      RECT 4.180000  0.285000 4.460000 0.615000 ;
      RECT 4.180000  0.615000 4.350000 0.715000 ;
      RECT 4.180000  0.885000 4.350000 1.825000 ;
      RECT 4.180000  1.995000 4.350000 2.065000 ;
      RECT 4.180000  2.065000 4.420000 2.440000 ;
      RECT 4.520000  0.780000 5.100000 1.035000 ;
      RECT 4.520000  1.035000 4.760000 1.905000 ;
      RECT 4.630000  0.705000 5.100000 0.780000 ;
      RECT 4.660000  2.190000 5.730000 2.360000 ;
      RECT 4.700000  0.365000 5.440000 0.535000 ;
      RECT 4.950000  1.655000 5.390000 2.010000 ;
      RECT 5.270000  0.535000 5.440000 1.315000 ;
      RECT 5.270000  1.315000 6.070000 1.485000 ;
      RECT 5.560000  1.485000 6.070000 1.575000 ;
      RECT 5.560000  1.575000 5.730000 2.190000 ;
      RECT 5.610000  0.765000 6.410000 1.065000 ;
      RECT 5.610000  1.065000 5.780000 1.095000 ;
      RECT 5.690000  0.085000 6.060000 0.585000 ;
      RECT 5.900000  1.245000 6.070000 1.315000 ;
      RECT 5.900000  1.835000 6.070000 2.635000 ;
      RECT 6.240000  0.365000 6.700000 0.535000 ;
      RECT 6.240000  0.535000 6.410000 0.765000 ;
      RECT 6.240000  1.065000 6.410000 2.135000 ;
      RECT 6.240000  2.135000 6.490000 2.465000 ;
      RECT 6.580000  0.705000 7.130000 1.035000 ;
      RECT 6.580000  1.245000 6.770000 1.965000 ;
      RECT 6.715000  2.165000 7.600000 2.335000 ;
      RECT 6.930000  0.365000 7.470000 0.535000 ;
      RECT 6.940000  1.035000 7.130000 1.575000 ;
      RECT 6.940000  1.575000 7.260000 1.905000 ;
      RECT 7.300000  0.535000 7.470000 0.995000 ;
      RECT 7.300000  0.995000 8.365000 1.325000 ;
      RECT 7.300000  1.325000 7.600000 1.405000 ;
      RECT 7.430000  1.405000 7.600000 2.165000 ;
      RECT 7.715000  0.085000 8.085000 0.615000 ;
      RECT 7.770000  1.575000 8.705000 1.905000 ;
      RECT 7.790000  2.135000 8.095000 2.635000 ;
      RECT 8.355000  0.300000 8.705000 0.825000 ;
      RECT 8.435000  1.905000 8.705000 2.455000 ;
      RECT 8.535000  0.825000 8.705000 0.995000 ;
      RECT 8.535000  0.995000 9.235000 1.325000 ;
      RECT 8.535000  1.325000 8.705000 1.575000 ;
      RECT 8.875000  0.085000 9.045000 0.695000 ;
      RECT 8.875000  1.625000 9.045000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.640000  1.785000 0.810000 1.955000 ;
      RECT 1.040000  0.765000 1.210000 0.935000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  0.765000 4.915000 0.935000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  1.785000 5.375000 1.955000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.590000  1.785000 6.760000 1.955000 ;
      RECT 6.630000  0.765000 6.800000 0.935000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 0.580000 1.755000 0.870000 1.800000 ;
      RECT 0.580000 1.800000 6.820000 1.940000 ;
      RECT 0.580000 1.940000 0.870000 1.985000 ;
      RECT 0.980000 0.735000 1.270000 0.780000 ;
      RECT 0.980000 0.780000 6.860000 0.920000 ;
      RECT 0.980000 0.920000 1.270000 0.965000 ;
      RECT 4.685000 0.735000 4.975000 0.780000 ;
      RECT 4.685000 0.920000 4.975000 0.965000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 6.530000 1.755000 6.820000 1.800000 ;
      RECT 6.530000 1.940000 6.820000 1.985000 ;
      RECT 6.570000 0.735000 6.860000 0.780000 ;
      RECT 6.570000 0.920000 6.860000 0.965000 ;
  END
END sky130_fd_sc_hd__sdfxtp_1
MACRO sky130_fd_sc_hd__sdfxtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.460000 1.355000 2.790000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.260000 0.305000 9.605000 0.820000 ;
        RECT 9.260000 1.505000 9.605000 2.395000 ;
        RECT 9.435000 0.820000 9.605000 1.505000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.530000 1.035000 4.020000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.780000 0.615000 3.250000 0.785000 ;
        RECT 1.780000 0.785000 1.950000 1.685000 ;
        RECT 2.475000 0.305000 2.650000 0.615000 ;
        RECT 3.080000 0.785000 3.250000 1.115000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.175000  0.345000  0.345000 0.635000 ;
      RECT 0.175000  0.635000  0.810000 0.805000 ;
      RECT 0.180000  1.795000  0.845000 1.965000 ;
      RECT 0.180000  1.965000  0.350000 2.465000 ;
      RECT 0.515000  0.085000  0.845000 0.465000 ;
      RECT 0.520000  2.135000  0.850000 2.635000 ;
      RECT 0.615000  0.805000  0.810000 0.970000 ;
      RECT 0.615000  0.970000  0.845000 1.795000 ;
      RECT 1.015000  0.345000  1.245000 0.715000 ;
      RECT 1.020000  0.715000  1.245000 2.465000 ;
      RECT 1.435000  0.275000  1.805000 0.445000 ;
      RECT 1.435000  0.445000  1.605000 1.860000 ;
      RECT 1.435000  1.860000  3.245000 2.075000 ;
      RECT 1.435000  2.075000  1.710000 2.445000 ;
      RECT 1.880000  2.245000  2.210000 2.635000 ;
      RECT 1.975000  0.085000  2.305000 0.445000 ;
      RECT 2.120000  0.955000  2.460000 1.125000 ;
      RECT 2.120000  1.125000  2.290000 1.860000 ;
      RECT 2.690000  2.245000  3.585000 2.415000 ;
      RECT 2.820000  0.275000  3.590000 0.445000 ;
      RECT 3.075000  1.355000  3.270000 1.685000 ;
      RECT 3.075000  1.685000  3.245000 1.860000 ;
      RECT 3.415000  1.825000  4.380000 1.995000 ;
      RECT 3.415000  1.995000  3.585000 2.245000 ;
      RECT 3.420000  0.445000  3.590000 0.695000 ;
      RECT 3.420000  0.695000  4.380000 0.865000 ;
      RECT 3.755000  2.165000  3.925000 2.635000 ;
      RECT 3.760000  0.085000  3.960000 0.525000 ;
      RECT 4.210000  0.365000  4.560000 0.535000 ;
      RECT 4.210000  0.535000  4.380000 0.695000 ;
      RECT 4.210000  0.865000  4.380000 1.825000 ;
      RECT 4.210000  1.995000  4.380000 2.065000 ;
      RECT 4.210000  2.065000  4.445000 2.440000 ;
      RECT 4.550000  0.705000  5.130000 1.035000 ;
      RECT 4.550000  1.035000  4.790000 1.905000 ;
      RECT 4.690000  2.190000  5.760000 2.360000 ;
      RECT 4.730000  0.365000  5.470000 0.535000 ;
      RECT 4.980000  1.655000  5.420000 2.010000 ;
      RECT 5.300000  0.535000  5.470000 1.315000 ;
      RECT 5.300000  1.315000  6.100000 1.485000 ;
      RECT 5.590000  1.485000  6.100000 1.575000 ;
      RECT 5.590000  1.575000  5.760000 2.190000 ;
      RECT 5.640000  0.765000  6.440000 1.065000 ;
      RECT 5.640000  1.065000  5.810000 1.095000 ;
      RECT 5.720000  0.085000  6.090000 0.585000 ;
      RECT 5.930000  1.245000  6.100000 1.315000 ;
      RECT 5.930000  1.835000  6.100000 2.635000 ;
      RECT 6.270000  0.365000  6.730000 0.535000 ;
      RECT 6.270000  0.535000  6.440000 0.765000 ;
      RECT 6.270000  1.065000  6.440000 2.135000 ;
      RECT 6.270000  2.135000  6.520000 2.465000 ;
      RECT 6.610000  0.705000  7.160000 1.035000 ;
      RECT 6.610000  1.245000  6.800000 1.965000 ;
      RECT 6.745000  2.165000  7.630000 2.335000 ;
      RECT 6.960000  0.365000  7.500000 0.535000 ;
      RECT 6.970000  1.035000  7.160000 1.575000 ;
      RECT 6.970000  1.575000  7.290000 1.905000 ;
      RECT 7.330000  0.535000  7.500000 0.995000 ;
      RECT 7.330000  0.995000  8.395000 1.325000 ;
      RECT 7.330000  1.325000  7.630000 1.405000 ;
      RECT 7.460000  1.405000  7.630000 2.165000 ;
      RECT 7.745000  0.085000  8.115000 0.615000 ;
      RECT 7.800000  1.575000  8.735000 1.905000 ;
      RECT 7.810000  2.135000  8.115000 2.635000 ;
      RECT 8.385000  0.300000  8.735000 0.825000 ;
      RECT 8.465000  1.905000  8.735000 2.455000 ;
      RECT 8.565000  0.825000  8.735000 0.995000 ;
      RECT 8.565000  0.995000  9.265000 1.325000 ;
      RECT 8.565000  1.325000  8.735000 1.575000 ;
      RECT 8.905000  0.085000  9.075000 0.695000 ;
      RECT 8.905000  1.625000  9.080000 2.635000 ;
      RECT 9.775000  0.085000  9.945000 0.930000 ;
      RECT 9.775000  1.405000  9.945000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.640000  1.785000 0.810000 1.955000 ;
      RECT 1.050000  0.765000 1.220000 0.935000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  0.765000 4.915000 0.935000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  1.785000 5.375000 1.955000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.620000  1.785000 6.790000 1.955000 ;
      RECT 6.630000  0.765000 6.800000 0.935000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
    LAYER met1 ;
      RECT 0.580000 1.755000 0.870000 1.800000 ;
      RECT 0.580000 1.800000 6.850000 1.940000 ;
      RECT 0.580000 1.940000 0.870000 1.985000 ;
      RECT 0.990000 0.735000 1.280000 0.780000 ;
      RECT 0.990000 0.780000 6.860000 0.920000 ;
      RECT 0.990000 0.920000 1.280000 0.965000 ;
      RECT 4.685000 0.735000 4.975000 0.780000 ;
      RECT 4.685000 0.920000 4.975000 0.965000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 6.560000 1.755000 6.850000 1.800000 ;
      RECT 6.560000 1.940000 6.850000 1.985000 ;
      RECT 6.570000 0.735000 6.860000 0.780000 ;
      RECT 6.570000 0.920000 6.860000 0.965000 ;
  END
END sky130_fd_sc_hd__sdfxtp_2
MACRO sky130_fd_sc_hd__sdfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.460000 1.355000 2.795000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.285000 0.305000  9.615000 0.735000 ;
        RECT  9.285000 0.735000 10.955000 0.905000 ;
        RECT  9.285000 1.505000 10.955000 1.675000 ;
        RECT  9.285000 1.675000  9.615000 2.395000 ;
        RECT 10.135000 0.305000 10.465000 0.735000 ;
        RECT 10.135000 1.675000 10.465000 2.395000 ;
        RECT 10.655000 0.905000 10.955000 1.505000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.535000 1.035000 4.025000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.780000 0.615000 3.255000 0.785000 ;
        RECT 1.780000 0.785000 1.950000 1.685000 ;
        RECT 2.475000 0.305000 2.650000 0.615000 ;
        RECT 3.085000 0.785000 3.255000 1.115000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.810000 0.805000 ;
      RECT  0.180000  1.795000  0.845000 1.965000 ;
      RECT  0.180000  1.965000  0.350000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.520000  2.135000  0.850000 2.635000 ;
      RECT  0.615000  0.805000  0.810000 0.970000 ;
      RECT  0.615000  0.970000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.245000 0.715000 ;
      RECT  1.020000  0.715000  1.245000 2.465000 ;
      RECT  1.435000  0.275000  1.805000 0.445000 ;
      RECT  1.435000  0.445000  1.605000 1.860000 ;
      RECT  1.435000  1.860000  3.250000 2.075000 ;
      RECT  1.435000  2.075000  1.710000 2.445000 ;
      RECT  1.880000  2.245000  2.210000 2.635000 ;
      RECT  1.975000  0.085000  2.305000 0.445000 ;
      RECT  2.120000  0.955000  2.465000 1.125000 ;
      RECT  2.120000  1.125000  2.290000 1.860000 ;
      RECT  2.695000  2.245000  3.590000 2.415000 ;
      RECT  2.820000  0.275000  3.595000 0.445000 ;
      RECT  3.080000  1.355000  3.275000 1.685000 ;
      RECT  3.080000  1.685000  3.250000 1.860000 ;
      RECT  3.420000  1.825000  4.385000 1.995000 ;
      RECT  3.420000  1.995000  3.590000 2.245000 ;
      RECT  3.425000  0.445000  3.595000 0.695000 ;
      RECT  3.425000  0.695000  4.385000 0.865000 ;
      RECT  3.760000  2.165000  3.930000 2.635000 ;
      RECT  3.765000  0.085000  3.965000 0.525000 ;
      RECT  4.215000  0.365000  4.565000 0.535000 ;
      RECT  4.215000  0.535000  4.385000 0.695000 ;
      RECT  4.215000  0.865000  4.385000 1.825000 ;
      RECT  4.215000  1.995000  4.385000 2.065000 ;
      RECT  4.215000  2.065000  4.450000 2.440000 ;
      RECT  4.555000  0.705000  5.135000 1.035000 ;
      RECT  4.555000  1.035000  4.795000 1.905000 ;
      RECT  4.695000  2.190000  5.765000 2.360000 ;
      RECT  4.735000  0.365000  5.475000 0.535000 ;
      RECT  4.985000  1.655000  5.425000 2.010000 ;
      RECT  5.305000  0.535000  5.475000 1.315000 ;
      RECT  5.305000  1.315000  6.105000 1.485000 ;
      RECT  5.595000  1.485000  6.105000 1.575000 ;
      RECT  5.595000  1.575000  5.765000 2.190000 ;
      RECT  5.645000  0.765000  6.445000 1.065000 ;
      RECT  5.645000  1.065000  5.815000 1.095000 ;
      RECT  5.725000  0.085000  6.095000 0.585000 ;
      RECT  5.935000  1.245000  6.105000 1.315000 ;
      RECT  5.935000  1.835000  6.105000 2.635000 ;
      RECT  6.275000  0.365000  6.735000 0.535000 ;
      RECT  6.275000  0.535000  6.445000 0.765000 ;
      RECT  6.275000  1.065000  6.445000 2.135000 ;
      RECT  6.275000  2.135000  6.525000 2.465000 ;
      RECT  6.615000  0.705000  7.165000 1.035000 ;
      RECT  6.615000  1.245000  6.805000 1.965000 ;
      RECT  6.750000  2.165000  7.635000 2.335000 ;
      RECT  6.965000  0.365000  7.505000 0.535000 ;
      RECT  6.975000  1.035000  7.165000 1.575000 ;
      RECT  6.975000  1.575000  7.295000 1.905000 ;
      RECT  7.335000  0.535000  7.505000 0.995000 ;
      RECT  7.335000  0.995000  8.400000 1.325000 ;
      RECT  7.335000  1.325000  7.635000 1.405000 ;
      RECT  7.465000  1.405000  7.635000 2.165000 ;
      RECT  7.750000  0.085000  8.120000 0.615000 ;
      RECT  7.805000  1.575000  8.755000 1.905000 ;
      RECT  7.815000  2.135000  8.120000 2.635000 ;
      RECT  8.390000  0.300000  8.750000 0.825000 ;
      RECT  8.470000  1.905000  8.755000 2.455000 ;
      RECT  8.570000  0.825000  8.750000 1.075000 ;
      RECT  8.570000  1.075000 10.485000 1.325000 ;
      RECT  8.570000  1.325000  8.755000 1.575000 ;
      RECT  8.925000  0.085000  9.095000 0.695000 ;
      RECT  8.925000  1.625000  9.105000 2.635000 ;
      RECT  9.795000  0.085000  9.965000 0.565000 ;
      RECT  9.795000  1.845000  9.965000 2.635000 ;
      RECT 10.635000  0.085000 10.805000 0.565000 ;
      RECT 10.635000  1.845000 10.805000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.615000  1.785000  0.785000 1.955000 ;
      RECT  1.055000  0.765000  1.225000 0.935000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.755000  0.765000  4.925000 0.935000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.215000  1.785000  5.385000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.625000  0.765000  6.795000 0.935000 ;
      RECT  6.625000  1.785000  6.795000 1.955000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 0.555000 1.755000 0.845000 1.800000 ;
      RECT 0.555000 1.800000 6.855000 1.940000 ;
      RECT 0.555000 1.940000 0.845000 1.985000 ;
      RECT 0.995000 0.735000 1.285000 0.780000 ;
      RECT 0.995000 0.780000 6.855000 0.920000 ;
      RECT 0.995000 0.920000 1.285000 0.965000 ;
      RECT 4.695000 0.735000 4.985000 0.780000 ;
      RECT 4.695000 0.920000 4.985000 0.965000 ;
      RECT 5.155000 1.755000 5.445000 1.800000 ;
      RECT 5.155000 1.940000 5.445000 1.985000 ;
      RECT 6.565000 0.735000 6.855000 0.780000 ;
      RECT 6.565000 0.920000 6.855000 0.965000 ;
      RECT 6.565000 1.755000 6.855000 1.800000 ;
      RECT 6.565000 1.940000 6.855000 1.985000 ;
  END
END sky130_fd_sc_hd__sdfxtp_4
MACRO sky130_fd_sc_hd__sdlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdlclkp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.850000 0.955000 1.190000 1.325000 ;
        RECT 0.880000 1.325000 1.190000 1.445000 ;
        RECT 0.880000 1.445000 1.235000 1.955000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.530000 0.255000 6.815000 0.825000 ;
        RECT 6.530000 1.495000 6.815000 2.465000 ;
        RECT 6.645000 0.825000 6.815000 1.495000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.340000 1.665000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.710000 0.955000 6.010000 1.265000 ;
        RECT 4.710000 1.265000 4.930000 1.325000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.090000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.615000 ;
      RECT 0.085000  0.615000 1.190000 0.785000 ;
      RECT 0.085000  1.835000 0.345000 2.635000 ;
      RECT 0.510000  0.785000 0.680000 1.460000 ;
      RECT 0.510000  1.460000 0.710000 1.755000 ;
      RECT 0.515000  0.085000 0.845000 0.445000 ;
      RECT 0.540000  1.755000 0.710000 2.125000 ;
      RECT 0.540000  2.125000 1.255000 2.465000 ;
      RECT 1.015000  0.255000 1.190000 0.615000 ;
      RECT 1.360000  0.255000 2.495000 0.535000 ;
      RECT 1.360000  0.705000 1.700000 1.205000 ;
      RECT 1.360000  1.205000 1.860000 1.325000 ;
      RECT 1.405000  1.325000 1.860000 1.955000 ;
      RECT 1.425000  2.125000 2.200000 2.465000 ;
      RECT 1.870000  0.705000 2.155000 1.035000 ;
      RECT 2.030000  1.205000 3.010000 1.375000 ;
      RECT 2.030000  1.375000 2.200000 2.125000 ;
      RECT 2.325000  0.535000 2.495000 0.995000 ;
      RECT 2.325000  0.995000 3.010000 1.205000 ;
      RECT 2.370000  1.575000 2.540000 1.635000 ;
      RECT 2.370000  1.635000 3.400000 1.905000 ;
      RECT 2.370000  2.075000 3.010000 2.635000 ;
      RECT 2.665000  0.085000 3.010000 0.825000 ;
      RECT 3.180000  0.255000 3.400000 1.635000 ;
      RECT 3.180000  1.905000 3.400000 1.915000 ;
      RECT 3.180000  1.915000 5.450000 2.085000 ;
      RECT 3.180000  2.085000 3.400000 2.465000 ;
      RECT 3.580000  0.255000 3.910000 0.765000 ;
      RECT 3.580000  0.765000 4.005000 0.935000 ;
      RECT 3.580000  0.935000 3.750000 1.575000 ;
      RECT 3.580000  1.575000 3.990000 1.745000 ;
      RECT 3.580000  2.255000 5.490000 2.635000 ;
      RECT 3.920000  1.105000 4.465000 1.275000 ;
      RECT 4.080000  0.085000 4.410000 0.445000 ;
      RECT 4.160000  1.275000 4.465000 1.495000 ;
      RECT 4.160000  1.495000 4.960000 1.745000 ;
      RECT 4.175000  0.615000 4.830000 0.785000 ;
      RECT 4.175000  0.785000 4.465000 1.105000 ;
      RECT 4.580000  0.255000 4.830000 0.615000 ;
      RECT 5.010000  0.255000 5.270000 0.615000 ;
      RECT 5.010000  0.615000 6.360000 0.785000 ;
      RECT 5.140000  1.435000 5.610000 1.605000 ;
      RECT 5.140000  1.605000 5.450000 1.915000 ;
      RECT 5.505000  0.085000 6.360000 0.445000 ;
      RECT 5.660000  1.775000 6.360000 2.085000 ;
      RECT 5.660000  2.085000 5.830000 2.465000 ;
      RECT 5.780000  1.435000 6.360000 1.775000 ;
      RECT 6.030000  2.255000 6.360000 2.635000 ;
      RECT 6.190000  0.785000 6.360000 0.995000 ;
      RECT 6.190000  0.995000 6.460000 1.325000 ;
      RECT 6.190000  1.325000 6.360000 1.435000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  1.445000 1.695000 1.615000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  0.765000 2.155000 0.935000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 3.835000  0.765000 4.005000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.295000  1.445000 4.465000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
    LAYER met1 ;
      RECT 1.465000 1.415000 1.755000 1.460000 ;
      RECT 1.465000 1.460000 4.525000 1.600000 ;
      RECT 1.465000 1.600000 1.755000 1.645000 ;
      RECT 1.925000 0.735000 2.215000 0.780000 ;
      RECT 1.925000 0.780000 4.065000 0.920000 ;
      RECT 1.925000 0.920000 2.215000 0.965000 ;
      RECT 3.775000 0.735000 4.065000 0.780000 ;
      RECT 3.775000 0.920000 4.065000 0.965000 ;
      RECT 4.235000 1.415000 4.525000 1.460000 ;
      RECT 4.235000 1.600000 4.525000 1.645000 ;
  END
END sky130_fd_sc_hd__sdlclkp_1
MACRO sky130_fd_sc_hd__sdlclkp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdlclkp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 0.955000 1.195000 1.445000 ;
        RECT 0.855000 1.445000 1.240000 1.955000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.570000 0.255000 6.840000 0.825000 ;
        RECT 6.570000 1.495000 6.840000 2.465000 ;
        RECT 6.670000 0.825000 6.840000 1.055000 ;
        RECT 6.670000 1.055000 7.275000 1.315000 ;
        RECT 6.670000 1.315000 6.840000 1.495000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.340000 1.665000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.705000 0.955000 6.050000 1.265000 ;
        RECT 4.705000 1.265000 4.925000 1.325000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.615000 ;
      RECT 0.085000  0.615000 1.195000 0.785000 ;
      RECT 0.085000  1.835000 0.345000 2.635000 ;
      RECT 0.515000  0.085000 0.845000 0.445000 ;
      RECT 0.515000  0.785000 0.685000 2.125000 ;
      RECT 0.515000  2.125000 1.260000 2.465000 ;
      RECT 1.015000  0.255000 1.195000 0.615000 ;
      RECT 1.365000  0.255000 2.500000 0.535000 ;
      RECT 1.365000  0.705000 1.705000 1.205000 ;
      RECT 1.365000  1.205000 1.865000 1.325000 ;
      RECT 1.410000  1.325000 1.865000 1.955000 ;
      RECT 1.430000  2.125000 2.205000 2.465000 ;
      RECT 1.875000  0.705000 2.160000 1.035000 ;
      RECT 2.035000  1.205000 3.015000 1.375000 ;
      RECT 2.035000  1.375000 2.205000 2.125000 ;
      RECT 2.330000  0.535000 2.500000 0.995000 ;
      RECT 2.330000  0.995000 3.015000 1.205000 ;
      RECT 2.375000  1.575000 2.545000 1.635000 ;
      RECT 2.375000  1.635000 3.405000 1.905000 ;
      RECT 2.375000  2.075000 3.015000 2.635000 ;
      RECT 2.670000  0.085000 3.015000 0.825000 ;
      RECT 3.185000  0.255000 3.405000 1.635000 ;
      RECT 3.185000  1.905000 3.405000 1.915000 ;
      RECT 3.185000  1.915000 5.490000 2.085000 ;
      RECT 3.185000  2.085000 3.405000 2.465000 ;
      RECT 3.575000  0.255000 3.925000 0.765000 ;
      RECT 3.575000  0.765000 4.000000 0.935000 ;
      RECT 3.575000  0.935000 3.745000 1.575000 ;
      RECT 3.575000  1.575000 4.040000 1.745000 ;
      RECT 3.575000  2.255000 5.530000 2.635000 ;
      RECT 3.915000  1.105000 4.460000 1.275000 ;
      RECT 4.095000  0.085000 4.425000 0.445000 ;
      RECT 4.170000  0.615000 4.825000 0.785000 ;
      RECT 4.170000  0.785000 4.460000 1.105000 ;
      RECT 4.210000  1.275000 4.460000 1.495000 ;
      RECT 4.210000  1.495000 5.010000 1.745000 ;
      RECT 4.595000  0.255000 4.825000 0.615000 ;
      RECT 5.100000  0.255000 5.310000 0.615000 ;
      RECT 5.100000  0.615000 6.400000 0.785000 ;
      RECT 5.180000  1.435000 5.650000 1.605000 ;
      RECT 5.180000  1.605000 5.490000 1.915000 ;
      RECT 5.490000  0.085000 6.400000 0.445000 ;
      RECT 5.700000  1.775000 6.400000 2.085000 ;
      RECT 5.700000  2.085000 5.870000 2.465000 ;
      RECT 5.820000  1.435000 6.400000 1.775000 ;
      RECT 6.070000  2.255000 6.400000 2.635000 ;
      RECT 6.230000  0.785000 6.400000 0.995000 ;
      RECT 6.230000  0.995000 6.500000 1.325000 ;
      RECT 6.230000  1.325000 6.400000 1.435000 ;
      RECT 7.010000  0.085000 7.275000 0.885000 ;
      RECT 7.010000  1.485000 7.275000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.530000  1.445000 1.700000 1.615000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 1.990000  0.765000 2.160000 0.935000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 3.830000  0.765000 4.000000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.290000  1.445000 4.460000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
    LAYER met1 ;
      RECT 1.470000 1.415000 1.760000 1.460000 ;
      RECT 1.470000 1.460000 4.520000 1.600000 ;
      RECT 1.470000 1.600000 1.760000 1.645000 ;
      RECT 1.930000 0.735000 2.220000 0.780000 ;
      RECT 1.930000 0.780000 4.060000 0.920000 ;
      RECT 1.930000 0.920000 2.220000 0.965000 ;
      RECT 3.770000 0.735000 4.060000 0.780000 ;
      RECT 3.770000 0.920000 4.060000 0.965000 ;
      RECT 4.230000 1.415000 4.520000 1.460000 ;
      RECT 4.230000 1.600000 4.520000 1.645000 ;
  END
END sky130_fd_sc_hd__sdlclkp_2
MACRO sky130_fd_sc_hd__sdlclkp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdlclkp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 0.955000 1.195000 1.445000 ;
        RECT 0.855000 1.445000 1.240000 1.955000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.500000 0.255000 6.830000 0.445000 ;
        RECT 6.580000 0.445000 6.830000 0.715000 ;
        RECT 6.580000 0.715000 7.220000 0.885000 ;
        RECT 6.580000 1.485000 7.220000 1.655000 ;
        RECT 6.580000 1.655000 6.830000 2.465000 ;
        RECT 7.050000 0.885000 7.220000 1.055000 ;
        RECT 7.050000 1.055000 8.195000 1.315000 ;
        RECT 7.050000 1.315000 7.220000 1.485000 ;
        RECT 7.420000 0.255000 7.720000 1.055000 ;
        RECT 7.420000 1.315000 7.720000 2.465000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.345000 1.665000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.406500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.725000 0.995000 4.945000 1.325000 ;
      LAYER mcon ;
        RECT 4.770000 1.105000 4.940000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.685000 0.995000 6.065000 1.325000 ;
      LAYER mcon ;
        RECT 5.710000 1.105000 5.880000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.710000 1.075000 5.000000 1.120000 ;
        RECT 4.710000 1.120000 5.940000 1.260000 ;
        RECT 4.710000 1.260000 5.000000 1.305000 ;
        RECT 5.650000 1.075000 5.940000 1.120000 ;
        RECT 5.650000 1.260000 5.940000 1.305000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.615000 ;
      RECT 0.085000  0.615000 1.195000 0.785000 ;
      RECT 0.085000  1.835000 0.345000 2.635000 ;
      RECT 0.515000  0.085000 0.845000 0.445000 ;
      RECT 0.515000  0.785000 0.685000 2.125000 ;
      RECT 0.515000  2.125000 1.260000 2.465000 ;
      RECT 1.015000  0.255000 1.195000 0.615000 ;
      RECT 1.365000  0.255000 2.500000 0.535000 ;
      RECT 1.365000  0.705000 1.705000 1.205000 ;
      RECT 1.365000  1.205000 1.865000 1.325000 ;
      RECT 1.410000  1.325000 1.865000 1.955000 ;
      RECT 1.430000  2.125000 2.205000 2.465000 ;
      RECT 1.875000  0.705000 2.160000 1.035000 ;
      RECT 2.035000  1.205000 3.015000 1.375000 ;
      RECT 2.035000  1.375000 2.205000 2.125000 ;
      RECT 2.330000  0.535000 2.500000 0.995000 ;
      RECT 2.330000  0.995000 3.015000 1.205000 ;
      RECT 2.375000  1.575000 2.545000 1.635000 ;
      RECT 2.375000  1.635000 3.405000 1.905000 ;
      RECT 2.375000  2.075000 3.015000 2.635000 ;
      RECT 2.670000  0.085000 3.015000 0.825000 ;
      RECT 3.185000  0.255000 3.405000 1.635000 ;
      RECT 3.185000  1.905000 3.405000 1.915000 ;
      RECT 3.185000  1.915000 5.515000 2.085000 ;
      RECT 3.185000  2.085000 3.405000 2.465000 ;
      RECT 3.595000  0.255000 3.925000 0.765000 ;
      RECT 3.595000  0.765000 4.020000 0.935000 ;
      RECT 3.595000  0.935000 3.765000 1.575000 ;
      RECT 3.595000  1.575000 4.005000 1.745000 ;
      RECT 3.595000  2.255000 5.515000 2.635000 ;
      RECT 3.935000  1.105000 4.480000 1.275000 ;
      RECT 4.095000  0.085000 4.425000 0.445000 ;
      RECT 4.175000  1.275000 4.480000 1.495000 ;
      RECT 4.175000  1.495000 4.975000 1.745000 ;
      RECT 4.190000  0.615000 4.845000 0.785000 ;
      RECT 4.190000  0.785000 4.480000 1.105000 ;
      RECT 4.595000  0.255000 4.845000 0.615000 ;
      RECT 5.015000  0.255000 5.435000 0.615000 ;
      RECT 5.015000  0.615000 6.410000 0.785000 ;
      RECT 5.165000  0.995000 5.515000 1.915000 ;
      RECT 5.605000  0.085000 6.330000 0.445000 ;
      RECT 5.685000  1.495000 6.410000 2.085000 ;
      RECT 5.685000  2.085000 5.855000 2.465000 ;
      RECT 6.055000  2.255000 6.385000 2.635000 ;
      RECT 6.240000  0.785000 6.410000 1.055000 ;
      RECT 6.240000  1.055000 6.880000 1.315000 ;
      RECT 6.240000  1.315000 6.410000 1.495000 ;
      RECT 7.000000  0.085000 7.250000 0.545000 ;
      RECT 7.000000  1.825000 7.250000 2.635000 ;
      RECT 7.890000  0.085000 8.195000 0.885000 ;
      RECT 7.890000  1.485000 8.195000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.530000  1.445000 1.700000 1.615000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 1.990000  0.765000 2.160000 0.935000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 3.850000  0.765000 4.020000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.310000  1.445000 4.480000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
    LAYER met1 ;
      RECT 1.470000 1.415000 1.760000 1.460000 ;
      RECT 1.470000 1.460000 4.540000 1.600000 ;
      RECT 1.470000 1.600000 1.760000 1.645000 ;
      RECT 1.930000 0.735000 2.220000 0.780000 ;
      RECT 1.930000 0.780000 4.080000 0.920000 ;
      RECT 1.930000 0.920000 2.220000 0.965000 ;
      RECT 3.790000 0.735000 4.080000 0.780000 ;
      RECT 3.790000 0.920000 4.080000 0.965000 ;
      RECT 4.250000 1.415000 4.540000 1.460000 ;
      RECT 4.250000 1.600000 4.540000 1.645000 ;
  END
END sky130_fd_sc_hd__sdlclkp_4
MACRO sky130_fd_sc_hd__sedfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.26000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.765000 1.915000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 0.765000 2.565000 1.185000 ;
        RECT 2.110000 1.185000 2.325000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.525000 0.255000 13.855000 2.420000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.700000 1.065000 12.145000 1.410000 ;
        RECT 11.700000 1.410000 12.030000 2.465000 ;
        RECT 11.815000 0.255000 12.145000 1.065000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 1.105000 6.215000 1.665000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025000 1.105000 5.250000 1.615000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.260000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  4.885000 1.435000 ;
        RECT -0.190000 1.435000 14.450000 2.910000 ;
        RECT  7.200000 1.305000 14.450000 1.435000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.260000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.260000 0.085000 ;
      RECT  0.000000  2.635000 14.260000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.845000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.355000  0.255000  1.785000 0.515000 ;
      RECT  1.355000  0.515000  1.525000 1.890000 ;
      RECT  1.355000  1.890000  1.785000 2.465000 ;
      RECT  2.235000  0.085000  2.565000 0.515000 ;
      RECT  2.235000  1.890000  2.565000 2.635000 ;
      RECT  2.495000  1.355000  3.085000 1.720000 ;
      RECT  2.755000  1.720000  3.085000 2.425000 ;
      RECT  2.780000  0.255000  3.005000 0.845000 ;
      RECT  2.780000  0.845000  3.635000 1.175000 ;
      RECT  2.780000  1.175000  3.085000 1.355000 ;
      RECT  3.185000  0.085000  3.515000 0.610000 ;
      RECT  3.265000  1.825000  3.460000 2.635000 ;
      RECT  3.805000  0.685000  3.975000 1.320000 ;
      RECT  3.805000  1.320000  4.175000 1.650000 ;
      RECT  4.125000  1.820000  4.515000 2.020000 ;
      RECT  4.125000  2.020000  4.455000 2.465000 ;
      RECT  4.145000  0.255000  4.415000 0.980000 ;
      RECT  4.145000  0.980000  4.515000 1.150000 ;
      RECT  4.345000  1.150000  4.515000 1.820000 ;
      RECT  4.595000  0.255000  4.795000 0.645000 ;
      RECT  4.595000  0.645000  4.855000 0.825000 ;
      RECT  4.635000  2.210000  4.965000 2.465000 ;
      RECT  4.685000  0.825000  4.855000 1.785000 ;
      RECT  4.685000  1.785000  4.965000 2.210000 ;
      RECT  4.965000  0.255000  5.590000 0.515000 ;
      RECT  5.155000  1.835000  6.585000 2.005000 ;
      RECT  5.155000  2.005000  5.495000 2.465000 ;
      RECT  5.260000  0.515000  5.590000 0.935000 ;
      RECT  5.420000  0.935000  5.590000 1.835000 ;
      RECT  5.665000  2.175000  6.010000 2.635000 ;
      RECT  5.760000  0.085000  6.010000 0.905000 ;
      RECT  6.385000  1.355000  6.585000 1.835000 ;
      RECT  6.515000  0.255000  7.135000 0.565000 ;
      RECT  6.515000  0.565000  6.925000 1.185000 ;
      RECT  6.675000  2.150000  7.005000 2.465000 ;
      RECT  6.755000  1.185000  6.925000 1.865000 ;
      RECT  6.755000  1.865000  7.005000 2.150000 ;
      RECT  7.095000  1.125000  7.280000 1.720000 ;
      RECT  7.115000  0.735000  7.620000 0.955000 ;
      RECT  7.215000  2.175000  8.255000 2.375000 ;
      RECT  7.305000  0.255000  7.980000 0.565000 ;
      RECT  7.450000  0.955000  7.620000 1.655000 ;
      RECT  7.450000  1.655000  7.915000 2.005000 ;
      RECT  7.810000  0.565000  7.980000 1.315000 ;
      RECT  7.810000  1.315000  8.660000 1.485000 ;
      RECT  8.085000  1.485000  8.660000 1.575000 ;
      RECT  8.085000  1.575000  8.255000 2.175000 ;
      RECT  8.170000  0.765000  9.235000 1.045000 ;
      RECT  8.170000  1.045000  9.745000 1.065000 ;
      RECT  8.170000  1.065000  8.370000 1.095000 ;
      RECT  8.245000  0.085000  8.640000 0.560000 ;
      RECT  8.425000  1.835000  8.660000 2.635000 ;
      RECT  8.490000  1.245000  8.660000 1.315000 ;
      RECT  8.830000  0.255000  9.235000 0.765000 ;
      RECT  8.830000  1.065000  9.745000 1.375000 ;
      RECT  8.830000  1.375000  9.160000 2.465000 ;
      RECT  9.370000  2.105000  9.660000 2.635000 ;
      RECT  9.465000  0.085000  9.740000 0.615000 ;
      RECT 10.090000  1.245000 10.280000 1.965000 ;
      RECT 10.225000  2.165000 11.190000 2.355000 ;
      RECT 10.305000  0.705000 10.770000 1.035000 ;
      RECT 10.325000  0.330000 11.190000 0.535000 ;
      RECT 10.450000  1.035000 10.770000 1.995000 ;
      RECT 10.940000  0.535000 11.190000 2.165000 ;
      RECT 11.360000  1.495000 11.530000 2.635000 ;
      RECT 11.395000  0.085000 11.645000 0.900000 ;
      RECT 12.200000  1.575000 12.430000 2.010000 ;
      RECT 12.315000  0.890000 12.940000 1.220000 ;
      RECT 12.600000  0.255000 12.940000 0.890000 ;
      RECT 12.600000  1.220000 12.940000 2.465000 ;
      RECT 13.110000  0.085000 13.355000 0.900000 ;
      RECT 13.110000  1.465000 13.355000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.635000  1.785000  0.805000 1.955000 ;
      RECT  1.015000  1.445000  1.185000 1.615000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.355000  0.425000  1.525000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.805000  0.765000  3.975000 0.935000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.185000  0.425000  4.355000 0.595000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.615000  0.425000  4.785000 0.595000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.530000  0.425000  6.700000 0.595000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.100000  1.445000  7.270000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.510000  1.785000  7.680000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.100000  1.785000 10.270000 1.955000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.520000  1.445000 10.690000 1.615000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 10.980000  1.785000 11.150000 1.955000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.230000  1.785000 12.400000 1.955000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 12.690000  0.765000 12.860000 0.935000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
    LAYER met1 ;
      RECT  0.575000 1.755000  0.865000 1.800000 ;
      RECT  0.575000 1.800000 10.330000 1.940000 ;
      RECT  0.575000 1.940000  0.865000 1.985000 ;
      RECT  0.955000 1.415000  1.245000 1.460000 ;
      RECT  0.955000 1.460000 10.750000 1.600000 ;
      RECT  0.955000 1.600000  1.245000 1.645000 ;
      RECT  1.295000 0.395000  4.415000 0.580000 ;
      RECT  1.295000 0.580000  1.585000 0.625000 ;
      RECT  3.745000 0.735000  4.035000 0.780000 ;
      RECT  3.745000 0.780000 12.920000 0.920000 ;
      RECT  3.745000 0.920000  4.035000 0.965000 ;
      RECT  4.125000 0.580000  4.415000 0.625000 ;
      RECT  4.555000 0.395000  6.760000 0.580000 ;
      RECT  4.555000 0.580000  4.845000 0.625000 ;
      RECT  6.470000 0.580000  6.760000 0.625000 ;
      RECT  7.040000 1.415000  7.330000 1.460000 ;
      RECT  7.040000 1.600000  7.330000 1.645000 ;
      RECT  7.450000 1.755000  7.740000 1.800000 ;
      RECT  7.450000 1.940000  7.740000 1.985000 ;
      RECT 10.040000 1.755000 10.330000 1.800000 ;
      RECT 10.040000 1.940000 10.330000 1.985000 ;
      RECT 10.460000 1.415000 10.750000 1.460000 ;
      RECT 10.460000 1.600000 10.750000 1.645000 ;
      RECT 10.920000 1.755000 11.210000 1.800000 ;
      RECT 10.920000 1.800000 12.460000 1.940000 ;
      RECT 10.920000 1.940000 11.210000 1.985000 ;
      RECT 12.170000 1.755000 12.460000 1.800000 ;
      RECT 12.170000 1.940000 12.460000 1.985000 ;
      RECT 12.630000 0.735000 12.920000 0.780000 ;
      RECT 12.630000 0.920000 12.920000 0.965000 ;
  END
END sky130_fd_sc_hd__sedfxbp_1
MACRO sky130_fd_sc_hd__sedfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.18000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.765000 1.915000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 0.765000 2.565000 1.185000 ;
        RECT 2.110000 1.185000 2.325000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.935000 0.255000 14.265000 2.420000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.700000 1.065000 12.145000 1.300000 ;
        RECT 11.700000 1.300000 12.030000 2.465000 ;
        RECT 11.815000 0.255000 12.145000 1.065000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 1.105000 6.215000 1.665000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025000 1.105000 5.250000 1.615000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 15.180000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  4.885000 1.435000 ;
        RECT -0.190000 1.435000 15.370000 2.910000 ;
        RECT  7.200000 1.305000 15.370000 1.435000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 15.180000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.180000 0.085000 ;
      RECT  0.000000  2.635000 15.180000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.845000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.355000  0.255000  1.785000 0.515000 ;
      RECT  1.355000  0.515000  1.525000 1.890000 ;
      RECT  1.355000  1.890000  1.785000 2.465000 ;
      RECT  2.235000  0.085000  2.565000 0.515000 ;
      RECT  2.235000  1.890000  2.565000 2.635000 ;
      RECT  2.495000  1.355000  3.085000 1.720000 ;
      RECT  2.755000  1.720000  3.085000 2.425000 ;
      RECT  2.780000  0.255000  3.005000 0.845000 ;
      RECT  2.780000  0.845000  3.635000 1.175000 ;
      RECT  2.780000  1.175000  3.085000 1.355000 ;
      RECT  3.185000  0.085000  3.515000 0.610000 ;
      RECT  3.265000  1.825000  3.460000 2.635000 ;
      RECT  3.805000  0.685000  3.975000 1.320000 ;
      RECT  3.805000  1.320000  4.175000 1.650000 ;
      RECT  4.125000  1.820000  4.515000 2.020000 ;
      RECT  4.125000  2.020000  4.455000 2.465000 ;
      RECT  4.145000  0.255000  4.415000 0.980000 ;
      RECT  4.145000  0.980000  4.515000 1.150000 ;
      RECT  4.345000  1.150000  4.515000 1.820000 ;
      RECT  4.595000  0.255000  4.795000 0.645000 ;
      RECT  4.595000  0.645000  4.855000 0.825000 ;
      RECT  4.635000  2.210000  4.965000 2.465000 ;
      RECT  4.685000  0.825000  4.855000 1.785000 ;
      RECT  4.685000  1.785000  4.965000 2.210000 ;
      RECT  4.965000  0.255000  5.590000 0.515000 ;
      RECT  5.155000  1.835000  6.585000 2.005000 ;
      RECT  5.155000  2.005000  5.495000 2.465000 ;
      RECT  5.260000  0.515000  5.590000 0.935000 ;
      RECT  5.420000  0.935000  5.590000 1.835000 ;
      RECT  5.665000  2.175000  6.010000 2.635000 ;
      RECT  5.760000  0.085000  6.010000 0.905000 ;
      RECT  6.385000  1.355000  6.585000 1.835000 ;
      RECT  6.515000  0.255000  7.135000 0.565000 ;
      RECT  6.515000  0.565000  6.925000 1.185000 ;
      RECT  6.675000  2.150000  7.005000 2.465000 ;
      RECT  6.755000  1.185000  6.925000 1.865000 ;
      RECT  6.755000  1.865000  7.005000 2.150000 ;
      RECT  7.095000  1.125000  7.280000 1.720000 ;
      RECT  7.115000  0.735000  7.620000 0.955000 ;
      RECT  7.215000  2.175000  8.255000 2.375000 ;
      RECT  7.305000  0.255000  7.980000 0.565000 ;
      RECT  7.450000  0.955000  7.620000 1.655000 ;
      RECT  7.450000  1.655000  7.915000 2.005000 ;
      RECT  7.810000  0.565000  7.980000 1.315000 ;
      RECT  7.810000  1.315000  8.660000 1.485000 ;
      RECT  8.085000  1.485000  8.660000 1.575000 ;
      RECT  8.085000  1.575000  8.255000 2.175000 ;
      RECT  8.170000  0.765000  9.235000 1.045000 ;
      RECT  8.170000  1.045000  9.745000 1.065000 ;
      RECT  8.170000  1.065000  8.370000 1.095000 ;
      RECT  8.245000  0.085000  8.640000 0.560000 ;
      RECT  8.425000  1.835000  8.660000 2.635000 ;
      RECT  8.490000  1.245000  8.660000 1.315000 ;
      RECT  8.830000  0.255000  9.235000 0.765000 ;
      RECT  8.830000  1.065000  9.745000 1.375000 ;
      RECT  8.830000  1.375000  9.160000 2.465000 ;
      RECT  9.370000  2.105000  9.660000 2.635000 ;
      RECT  9.465000  0.085000  9.740000 0.615000 ;
      RECT 10.090000  1.245000 10.280000 1.965000 ;
      RECT 10.225000  2.165000 11.190000 2.355000 ;
      RECT 10.305000  0.705000 10.770000 1.035000 ;
      RECT 10.325000  0.330000 11.190000 0.535000 ;
      RECT 10.450000  1.035000 10.770000 1.995000 ;
      RECT 10.940000  0.535000 11.190000 2.165000 ;
      RECT 11.360000  1.495000 11.530000 2.635000 ;
      RECT 11.395000  0.085000 11.645000 0.900000 ;
      RECT 12.200000  1.465000 12.450000 2.635000 ;
      RECT 12.315000  0.085000 12.565000 0.900000 ;
      RECT 12.620000  1.575000 12.850000 2.010000 ;
      RECT 12.735000  0.890000 13.360000 1.220000 ;
      RECT 13.020000  0.255000 13.360000 0.890000 ;
      RECT 13.020000  1.220000 13.360000 2.465000 ;
      RECT 13.530000  0.085000 13.765000 0.900000 ;
      RECT 13.530000  1.465000 13.765000 2.635000 ;
      RECT 14.435000  0.085000 14.695000 0.900000 ;
      RECT 14.435000  1.465000 14.695000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.635000  1.785000  0.805000 1.955000 ;
      RECT  1.015000  1.445000  1.185000 1.615000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.355000  0.425000  1.525000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.805000  0.765000  3.975000 0.935000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.185000  0.425000  4.355000 0.595000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.615000  0.425000  4.785000 0.595000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.530000  0.425000  6.700000 0.595000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.100000  1.445000  7.270000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.510000  1.785000  7.680000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.100000  1.785000 10.270000 1.955000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.520000  1.445000 10.690000 1.615000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 10.980000  1.785000 11.150000 1.955000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 12.650000  1.785000 12.820000 1.955000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.110000  0.765000 13.280000 0.935000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
    LAYER met1 ;
      RECT  0.575000 1.755000  0.865000 1.800000 ;
      RECT  0.575000 1.800000 10.330000 1.940000 ;
      RECT  0.575000 1.940000  0.865000 1.985000 ;
      RECT  0.955000 1.415000  1.245000 1.460000 ;
      RECT  0.955000 1.460000 10.750000 1.600000 ;
      RECT  0.955000 1.600000  1.245000 1.645000 ;
      RECT  1.295000 0.395000  4.415000 0.580000 ;
      RECT  1.295000 0.580000  1.585000 0.625000 ;
      RECT  3.745000 0.735000  4.035000 0.780000 ;
      RECT  3.745000 0.780000 13.340000 0.920000 ;
      RECT  3.745000 0.920000  4.035000 0.965000 ;
      RECT  4.125000 0.580000  4.415000 0.625000 ;
      RECT  4.555000 0.395000  6.760000 0.580000 ;
      RECT  4.555000 0.580000  4.845000 0.625000 ;
      RECT  6.470000 0.580000  6.760000 0.625000 ;
      RECT  7.040000 1.415000  7.330000 1.460000 ;
      RECT  7.040000 1.600000  7.330000 1.645000 ;
      RECT  7.450000 1.755000  7.740000 1.800000 ;
      RECT  7.450000 1.940000  7.740000 1.985000 ;
      RECT 10.040000 1.755000 10.330000 1.800000 ;
      RECT 10.040000 1.940000 10.330000 1.985000 ;
      RECT 10.460000 1.415000 10.750000 1.460000 ;
      RECT 10.460000 1.600000 10.750000 1.645000 ;
      RECT 10.920000 1.755000 11.210000 1.800000 ;
      RECT 10.920000 1.800000 12.880000 1.940000 ;
      RECT 10.920000 1.940000 11.210000 1.985000 ;
      RECT 12.590000 1.755000 12.880000 1.800000 ;
      RECT 12.590000 1.940000 12.880000 1.985000 ;
      RECT 13.050000 0.735000 13.340000 0.780000 ;
      RECT 13.050000 0.920000 13.340000 0.965000 ;
  END
END sky130_fd_sc_hd__sedfxbp_2
MACRO sky130_fd_sc_hd__sedfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.34000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.765000 1.915000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 0.765000 2.565000 1.185000 ;
        RECT 2.110000 1.185000 2.325000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.765000 0.305000 13.095000 2.420000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 1.105000 6.215000 1.665000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025000 1.105000 5.250000 1.615000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.340000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  4.885000 1.435000 ;
        RECT -0.190000 1.435000 13.530000 2.910000 ;
        RECT  7.200000 1.305000 13.530000 1.435000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.340000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.340000 0.085000 ;
      RECT  0.000000  2.635000 13.340000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.845000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.355000  0.255000  1.785000 0.515000 ;
      RECT  1.355000  0.515000  1.525000 1.890000 ;
      RECT  1.355000  1.890000  1.785000 2.465000 ;
      RECT  2.235000  0.085000  2.565000 0.515000 ;
      RECT  2.235000  1.890000  2.565000 2.635000 ;
      RECT  2.495000  1.355000  3.085000 1.720000 ;
      RECT  2.755000  1.720000  3.085000 2.425000 ;
      RECT  2.780000  0.255000  3.005000 0.845000 ;
      RECT  2.780000  0.845000  3.635000 1.175000 ;
      RECT  2.780000  1.175000  3.085000 1.355000 ;
      RECT  3.185000  0.085000  3.515000 0.610000 ;
      RECT  3.265000  1.825000  3.460000 2.635000 ;
      RECT  3.805000  0.685000  3.975000 1.320000 ;
      RECT  3.805000  1.320000  4.175000 1.650000 ;
      RECT  4.125000  1.820000  4.515000 2.020000 ;
      RECT  4.125000  2.020000  4.455000 2.465000 ;
      RECT  4.145000  0.255000  4.415000 0.980000 ;
      RECT  4.145000  0.980000  4.515000 1.150000 ;
      RECT  4.345000  1.150000  4.515000 1.820000 ;
      RECT  4.595000  0.255000  4.795000 0.645000 ;
      RECT  4.595000  0.645000  4.855000 0.825000 ;
      RECT  4.635000  2.210000  4.965000 2.465000 ;
      RECT  4.685000  0.825000  4.855000 1.785000 ;
      RECT  4.685000  1.785000  4.965000 2.210000 ;
      RECT  4.965000  0.255000  5.590000 0.515000 ;
      RECT  5.155000  1.835000  6.585000 2.005000 ;
      RECT  5.155000  2.005000  5.495000 2.465000 ;
      RECT  5.260000  0.515000  5.590000 0.935000 ;
      RECT  5.420000  0.935000  5.590000 1.835000 ;
      RECT  5.665000  2.175000  6.010000 2.635000 ;
      RECT  5.760000  0.085000  6.010000 0.905000 ;
      RECT  6.385000  1.355000  6.585000 1.835000 ;
      RECT  6.515000  0.255000  7.135000 0.565000 ;
      RECT  6.515000  0.565000  6.925000 1.185000 ;
      RECT  6.675000  2.150000  7.005000 2.465000 ;
      RECT  6.755000  1.185000  6.925000 1.865000 ;
      RECT  6.755000  1.865000  7.005000 2.150000 ;
      RECT  7.095000  1.125000  7.280000 1.720000 ;
      RECT  7.115000  0.735000  7.620000 0.955000 ;
      RECT  7.215000  2.175000  8.255000 2.375000 ;
      RECT  7.305000  0.255000  7.980000 0.565000 ;
      RECT  7.450000  0.955000  7.620000 1.655000 ;
      RECT  7.450000  1.655000  7.915000 2.005000 ;
      RECT  7.810000  0.565000  7.980000 1.315000 ;
      RECT  7.810000  1.315000  8.660000 1.485000 ;
      RECT  8.085000  1.485000  8.660000 1.575000 ;
      RECT  8.085000  1.575000  8.255000 2.175000 ;
      RECT  8.170000  0.765000  9.235000 1.045000 ;
      RECT  8.170000  1.045000  9.745000 1.065000 ;
      RECT  8.170000  1.065000  8.370000 1.095000 ;
      RECT  8.245000  0.085000  8.640000 0.560000 ;
      RECT  8.425000  1.835000  8.660000 2.635000 ;
      RECT  8.490000  1.245000  8.660000 1.315000 ;
      RECT  8.830000  0.255000  9.235000 0.765000 ;
      RECT  8.830000  1.065000  9.745000 1.375000 ;
      RECT  8.830000  1.375000  9.160000 2.465000 ;
      RECT  9.370000  2.105000  9.660000 2.635000 ;
      RECT  9.465000  0.085000  9.740000 0.615000 ;
      RECT 10.090000  1.245000 10.280000 1.965000 ;
      RECT 10.225000  2.165000 11.110000 2.355000 ;
      RECT 10.305000  0.705000 10.770000 1.035000 ;
      RECT 10.325000  0.330000 11.110000 0.535000 ;
      RECT 10.450000  1.035000 10.770000 1.995000 ;
      RECT 10.940000  0.535000 11.110000 0.995000 ;
      RECT 10.940000  0.995000 11.810000 1.325000 ;
      RECT 10.940000  1.325000 11.110000 2.165000 ;
      RECT 11.280000  1.530000 12.180000 1.905000 ;
      RECT 11.280000  2.135000 11.540000 2.635000 ;
      RECT 11.350000  0.085000 11.665000 0.615000 ;
      RECT 11.840000  1.905000 12.180000 2.465000 ;
      RECT 11.850000  0.300000 12.180000 0.825000 ;
      RECT 11.990000  0.825000 12.180000 1.530000 ;
      RECT 12.350000  0.085000 12.595000 0.900000 ;
      RECT 12.350000  1.465000 12.595000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.635000  1.785000  0.805000 1.955000 ;
      RECT  1.015000  1.445000  1.185000 1.615000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.355000  0.425000  1.525000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.805000  0.765000  3.975000 0.935000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.185000  0.425000  4.355000 0.595000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.615000  0.425000  4.785000 0.595000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.530000  0.425000  6.700000 0.595000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.100000  1.445000  7.270000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.510000  1.785000  7.680000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.100000  1.785000 10.270000 1.955000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.520000  1.445000 10.690000 1.615000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.000000  0.765000 12.170000 0.935000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
    LAYER met1 ;
      RECT  0.575000 1.755000  0.865000 1.800000 ;
      RECT  0.575000 1.800000 10.330000 1.940000 ;
      RECT  0.575000 1.940000  0.865000 1.985000 ;
      RECT  0.955000 1.415000  1.245000 1.460000 ;
      RECT  0.955000 1.460000 10.750000 1.600000 ;
      RECT  0.955000 1.600000  1.245000 1.645000 ;
      RECT  1.295000 0.395000  4.415000 0.580000 ;
      RECT  1.295000 0.580000  1.585000 0.625000 ;
      RECT  3.745000 0.735000  4.035000 0.780000 ;
      RECT  3.745000 0.780000 12.230000 0.920000 ;
      RECT  3.745000 0.920000  4.035000 0.965000 ;
      RECT  4.125000 0.580000  4.415000 0.625000 ;
      RECT  4.555000 0.395000  6.760000 0.580000 ;
      RECT  4.555000 0.580000  4.845000 0.625000 ;
      RECT  6.470000 0.580000  6.760000 0.625000 ;
      RECT  7.040000 1.415000  7.330000 1.460000 ;
      RECT  7.040000 1.600000  7.330000 1.645000 ;
      RECT  7.450000 1.755000  7.740000 1.800000 ;
      RECT  7.450000 1.940000  7.740000 1.985000 ;
      RECT 10.040000 1.755000 10.330000 1.800000 ;
      RECT 10.040000 1.940000 10.330000 1.985000 ;
      RECT 10.460000 1.415000 10.750000 1.460000 ;
      RECT 10.460000 1.600000 10.750000 1.645000 ;
      RECT 11.940000 0.735000 12.230000 0.780000 ;
      RECT 11.940000 0.920000 12.230000 0.965000 ;
  END
END sky130_fd_sc_hd__sedfxtp_1
MACRO sky130_fd_sc_hd__sedfxtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.80000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.765000 1.915000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 0.765000 2.565000 1.185000 ;
        RECT 2.110000 1.185000 2.325000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.755000 0.305000 13.085000 2.420000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 1.105000 6.215000 1.665000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025000 1.105000 5.250000 1.615000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.800000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  4.885000 1.435000 ;
        RECT -0.190000 1.435000 13.990000 2.910000 ;
        RECT  7.200000 1.305000 13.990000 1.435000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.800000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.800000 0.085000 ;
      RECT  0.000000  2.635000 13.800000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.845000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.355000  0.255000  1.785000 0.515000 ;
      RECT  1.355000  0.515000  1.525000 1.890000 ;
      RECT  1.355000  1.890000  1.785000 2.465000 ;
      RECT  2.235000  0.085000  2.565000 0.515000 ;
      RECT  2.235000  1.890000  2.565000 2.635000 ;
      RECT  2.495000  1.355000  3.085000 1.720000 ;
      RECT  2.755000  1.720000  3.085000 2.425000 ;
      RECT  2.780000  0.255000  3.005000 0.845000 ;
      RECT  2.780000  0.845000  3.635000 1.175000 ;
      RECT  2.780000  1.175000  3.085000 1.355000 ;
      RECT  3.185000  0.085000  3.515000 0.610000 ;
      RECT  3.265000  1.825000  3.460000 2.635000 ;
      RECT  3.805000  0.685000  3.975000 1.320000 ;
      RECT  3.805000  1.320000  4.175000 1.650000 ;
      RECT  4.125000  1.820000  4.515000 2.020000 ;
      RECT  4.125000  2.020000  4.455000 2.465000 ;
      RECT  4.145000  0.255000  4.415000 0.980000 ;
      RECT  4.145000  0.980000  4.515000 1.150000 ;
      RECT  4.345000  1.150000  4.515000 1.820000 ;
      RECT  4.595000  0.255000  4.795000 0.645000 ;
      RECT  4.595000  0.645000  4.855000 0.825000 ;
      RECT  4.635000  2.210000  4.965000 2.465000 ;
      RECT  4.685000  0.825000  4.855000 1.785000 ;
      RECT  4.685000  1.785000  4.965000 2.210000 ;
      RECT  4.965000  0.255000  5.590000 0.515000 ;
      RECT  5.155000  1.835000  6.585000 2.005000 ;
      RECT  5.155000  2.005000  5.495000 2.465000 ;
      RECT  5.260000  0.515000  5.590000 0.935000 ;
      RECT  5.420000  0.935000  5.590000 1.835000 ;
      RECT  5.665000  2.175000  6.010000 2.635000 ;
      RECT  5.760000  0.085000  6.010000 0.905000 ;
      RECT  6.385000  1.355000  6.585000 1.835000 ;
      RECT  6.515000  0.255000  7.135000 0.565000 ;
      RECT  6.515000  0.565000  6.925000 1.185000 ;
      RECT  6.675000  2.150000  7.005000 2.465000 ;
      RECT  6.755000  1.185000  6.925000 1.865000 ;
      RECT  6.755000  1.865000  7.005000 2.150000 ;
      RECT  7.095000  1.125000  7.280000 1.720000 ;
      RECT  7.115000  0.735000  7.620000 0.955000 ;
      RECT  7.215000  2.175000  8.255000 2.375000 ;
      RECT  7.305000  0.255000  7.980000 0.565000 ;
      RECT  7.450000  0.955000  7.620000 1.655000 ;
      RECT  7.450000  1.655000  7.915000 2.005000 ;
      RECT  7.810000  0.565000  7.980000 1.315000 ;
      RECT  7.810000  1.315000  8.660000 1.485000 ;
      RECT  8.085000  1.485000  8.660000 1.575000 ;
      RECT  8.085000  1.575000  8.255000 2.175000 ;
      RECT  8.170000  0.765000  9.235000 1.045000 ;
      RECT  8.170000  1.045000  9.745000 1.065000 ;
      RECT  8.170000  1.065000  8.370000 1.095000 ;
      RECT  8.245000  0.085000  8.640000 0.560000 ;
      RECT  8.425000  1.835000  8.660000 2.635000 ;
      RECT  8.490000  1.245000  8.660000 1.315000 ;
      RECT  8.830000  0.255000  9.235000 0.765000 ;
      RECT  8.830000  1.065000  9.745000 1.375000 ;
      RECT  8.830000  1.375000  9.160000 2.465000 ;
      RECT  9.370000  2.105000  9.660000 2.635000 ;
      RECT  9.465000  0.085000  9.740000 0.615000 ;
      RECT 10.090000  1.245000 10.280000 1.965000 ;
      RECT 10.225000  2.165000 11.110000 2.355000 ;
      RECT 10.305000  0.705000 10.770000 1.035000 ;
      RECT 10.325000  0.330000 11.110000 0.535000 ;
      RECT 10.450000  1.035000 10.770000 1.995000 ;
      RECT 10.940000  0.535000 11.110000 0.995000 ;
      RECT 10.940000  0.995000 11.810000 1.325000 ;
      RECT 10.940000  1.325000 11.110000 2.165000 ;
      RECT 11.280000  1.530000 12.180000 1.905000 ;
      RECT 11.280000  2.135000 11.540000 2.635000 ;
      RECT 11.350000  0.085000 11.665000 0.615000 ;
      RECT 11.840000  1.905000 12.180000 2.465000 ;
      RECT 11.850000  0.300000 12.180000 0.825000 ;
      RECT 11.990000  0.825000 12.180000 1.530000 ;
      RECT 12.350000  0.085000 12.585000 0.900000 ;
      RECT 12.350000  1.465000 12.585000 2.635000 ;
      RECT 13.255000  0.085000 13.515000 0.900000 ;
      RECT 13.255000  1.465000 13.515000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.635000  1.785000  0.805000 1.955000 ;
      RECT  1.015000  1.445000  1.185000 1.615000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.355000  0.425000  1.525000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.805000  0.765000  3.975000 0.935000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.185000  0.425000  4.355000 0.595000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.615000  0.425000  4.785000 0.595000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.530000  0.425000  6.700000 0.595000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.100000  1.445000  7.270000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.510000  1.785000  7.680000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.100000  1.785000 10.270000 1.955000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.520000  1.445000 10.690000 1.615000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.000000  0.765000 12.170000 0.935000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
    LAYER met1 ;
      RECT  0.575000 1.755000  0.865000 1.800000 ;
      RECT  0.575000 1.800000 10.330000 1.940000 ;
      RECT  0.575000 1.940000  0.865000 1.985000 ;
      RECT  0.955000 1.415000  1.245000 1.460000 ;
      RECT  0.955000 1.460000 10.750000 1.600000 ;
      RECT  0.955000 1.600000  1.245000 1.645000 ;
      RECT  1.295000 0.395000  4.415000 0.580000 ;
      RECT  1.295000 0.580000  1.585000 0.625000 ;
      RECT  3.745000 0.735000  4.035000 0.780000 ;
      RECT  3.745000 0.780000 12.230000 0.920000 ;
      RECT  3.745000 0.920000  4.035000 0.965000 ;
      RECT  4.125000 0.580000  4.415000 0.625000 ;
      RECT  4.555000 0.395000  6.760000 0.580000 ;
      RECT  4.555000 0.580000  4.845000 0.625000 ;
      RECT  6.470000 0.580000  6.760000 0.625000 ;
      RECT  7.040000 1.415000  7.330000 1.460000 ;
      RECT  7.040000 1.600000  7.330000 1.645000 ;
      RECT  7.450000 1.755000  7.740000 1.800000 ;
      RECT  7.450000 1.940000  7.740000 1.985000 ;
      RECT 10.040000 1.755000 10.330000 1.800000 ;
      RECT 10.040000 1.940000 10.330000 1.985000 ;
      RECT 10.460000 1.415000 10.750000 1.460000 ;
      RECT 10.460000 1.600000 10.750000 1.645000 ;
      RECT 11.940000 0.735000 12.230000 0.780000 ;
      RECT 11.940000 0.920000 12.230000 0.965000 ;
  END
END sky130_fd_sc_hd__sedfxtp_2
MACRO sky130_fd_sc_hd__sedfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.72000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.765000 1.915000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 0.765000 2.565000 1.185000 ;
        RECT 2.110000 1.185000 2.325000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.755000 0.305000 13.085000 1.070000 ;
        RECT 12.755000 1.070000 13.925000 1.295000 ;
        RECT 12.755000 1.295000 13.085000 2.420000 ;
        RECT 13.595000 0.305000 13.925000 1.070000 ;
        RECT 13.595000 1.295000 13.925000 2.420000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 1.105000 6.215000 1.665000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025000 1.105000 5.250000 1.615000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.720000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  4.885000 1.435000 ;
        RECT -0.190000 1.435000 14.910000 2.910000 ;
        RECT  7.200000 1.305000 14.910000 1.435000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.720000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.720000 0.085000 ;
      RECT  0.000000  2.635000 14.720000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.845000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.355000  0.255000  1.785000 0.515000 ;
      RECT  1.355000  0.515000  1.525000 1.890000 ;
      RECT  1.355000  1.890000  1.785000 2.465000 ;
      RECT  2.235000  0.085000  2.565000 0.515000 ;
      RECT  2.235000  1.890000  2.565000 2.635000 ;
      RECT  2.495000  1.355000  3.085000 1.720000 ;
      RECT  2.755000  1.720000  3.085000 2.425000 ;
      RECT  2.780000  0.255000  3.005000 0.845000 ;
      RECT  2.780000  0.845000  3.635000 1.175000 ;
      RECT  2.780000  1.175000  3.085000 1.355000 ;
      RECT  3.185000  0.085000  3.515000 0.610000 ;
      RECT  3.265000  1.825000  3.460000 2.635000 ;
      RECT  3.805000  0.685000  3.975000 1.320000 ;
      RECT  3.805000  1.320000  4.175000 1.650000 ;
      RECT  4.125000  1.820000  4.515000 2.020000 ;
      RECT  4.125000  2.020000  4.455000 2.465000 ;
      RECT  4.145000  0.255000  4.415000 0.980000 ;
      RECT  4.145000  0.980000  4.515000 1.150000 ;
      RECT  4.345000  1.150000  4.515000 1.820000 ;
      RECT  4.595000  0.255000  4.795000 0.645000 ;
      RECT  4.595000  0.645000  4.855000 0.825000 ;
      RECT  4.635000  2.210000  4.965000 2.465000 ;
      RECT  4.685000  0.825000  4.855000 1.785000 ;
      RECT  4.685000  1.785000  4.965000 2.210000 ;
      RECT  4.965000  0.255000  5.590000 0.515000 ;
      RECT  5.155000  1.835000  6.585000 2.005000 ;
      RECT  5.155000  2.005000  5.495000 2.465000 ;
      RECT  5.260000  0.515000  5.590000 0.935000 ;
      RECT  5.420000  0.935000  5.590000 1.835000 ;
      RECT  5.665000  2.175000  6.010000 2.635000 ;
      RECT  5.760000  0.085000  6.010000 0.905000 ;
      RECT  6.385000  1.355000  6.585000 1.835000 ;
      RECT  6.515000  0.255000  7.135000 0.565000 ;
      RECT  6.515000  0.565000  6.925000 1.185000 ;
      RECT  6.675000  2.150000  7.005000 2.465000 ;
      RECT  6.755000  1.185000  6.925000 1.865000 ;
      RECT  6.755000  1.865000  7.005000 2.150000 ;
      RECT  7.095000  1.125000  7.280000 1.720000 ;
      RECT  7.115000  0.735000  7.620000 0.955000 ;
      RECT  7.215000  2.175000  8.255000 2.375000 ;
      RECT  7.305000  0.255000  7.980000 0.565000 ;
      RECT  7.450000  0.955000  7.620000 1.655000 ;
      RECT  7.450000  1.655000  7.915000 2.005000 ;
      RECT  7.810000  0.565000  7.980000 1.315000 ;
      RECT  7.810000  1.315000  8.660000 1.485000 ;
      RECT  8.085000  1.485000  8.660000 1.575000 ;
      RECT  8.085000  1.575000  8.255000 2.175000 ;
      RECT  8.170000  0.765000  9.235000 1.045000 ;
      RECT  8.170000  1.045000  9.745000 1.065000 ;
      RECT  8.170000  1.065000  8.370000 1.095000 ;
      RECT  8.245000  0.085000  8.640000 0.560000 ;
      RECT  8.425000  1.835000  8.660000 2.635000 ;
      RECT  8.490000  1.245000  8.660000 1.315000 ;
      RECT  8.830000  0.255000  9.235000 0.765000 ;
      RECT  8.830000  1.065000  9.745000 1.375000 ;
      RECT  8.830000  1.375000  9.160000 2.465000 ;
      RECT  9.370000  2.105000  9.660000 2.635000 ;
      RECT  9.465000  0.085000  9.740000 0.615000 ;
      RECT 10.090000  1.245000 10.280000 1.965000 ;
      RECT 10.225000  2.165000 11.110000 2.355000 ;
      RECT 10.305000  0.705000 10.770000 1.035000 ;
      RECT 10.325000  0.330000 11.110000 0.535000 ;
      RECT 10.450000  1.035000 10.770000 1.995000 ;
      RECT 10.940000  0.535000 11.110000 0.995000 ;
      RECT 10.940000  0.995000 11.810000 1.325000 ;
      RECT 10.940000  1.325000 11.110000 2.165000 ;
      RECT 11.280000  1.530000 12.180000 1.905000 ;
      RECT 11.280000  2.135000 11.540000 2.635000 ;
      RECT 11.350000  0.085000 11.665000 0.615000 ;
      RECT 11.840000  1.905000 12.180000 2.465000 ;
      RECT 11.850000  0.300000 12.180000 0.825000 ;
      RECT 11.990000  0.825000 12.180000 1.530000 ;
      RECT 12.350000  0.085000 12.585000 0.900000 ;
      RECT 12.350000  1.465000 12.585000 2.635000 ;
      RECT 13.255000  0.085000 13.425000 0.900000 ;
      RECT 13.255000  1.465000 13.425000 2.635000 ;
      RECT 14.095000  0.085000 14.355000 1.280000 ;
      RECT 14.095000  1.465000 14.355000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.635000  1.785000  0.805000 1.955000 ;
      RECT  1.015000  1.445000  1.185000 1.615000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.355000  0.425000  1.525000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.805000  0.765000  3.975000 0.935000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.185000  0.425000  4.355000 0.595000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.615000  0.425000  4.785000 0.595000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.530000  0.425000  6.700000 0.595000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.100000  1.445000  7.270000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.510000  1.785000  7.680000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.100000  1.785000 10.270000 1.955000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.520000  1.445000 10.690000 1.615000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.000000  0.765000 12.170000 0.935000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
    LAYER met1 ;
      RECT  0.575000 1.755000  0.865000 1.800000 ;
      RECT  0.575000 1.800000 10.330000 1.940000 ;
      RECT  0.575000 1.940000  0.865000 1.985000 ;
      RECT  0.955000 1.415000  1.245000 1.460000 ;
      RECT  0.955000 1.460000 10.750000 1.600000 ;
      RECT  0.955000 1.600000  1.245000 1.645000 ;
      RECT  1.295000 0.395000  4.415000 0.580000 ;
      RECT  1.295000 0.580000  1.585000 0.625000 ;
      RECT  3.745000 0.735000  4.035000 0.780000 ;
      RECT  3.745000 0.780000 12.230000 0.920000 ;
      RECT  3.745000 0.920000  4.035000 0.965000 ;
      RECT  4.125000 0.580000  4.415000 0.625000 ;
      RECT  4.555000 0.395000  6.760000 0.580000 ;
      RECT  4.555000 0.580000  4.845000 0.625000 ;
      RECT  6.470000 0.580000  6.760000 0.625000 ;
      RECT  7.040000 1.415000  7.330000 1.460000 ;
      RECT  7.040000 1.600000  7.330000 1.645000 ;
      RECT  7.450000 1.755000  7.740000 1.800000 ;
      RECT  7.450000 1.940000  7.740000 1.985000 ;
      RECT 10.040000 1.755000 10.330000 1.800000 ;
      RECT 10.040000 1.940000 10.330000 1.985000 ;
      RECT 10.460000 1.415000 10.750000 1.460000 ;
      RECT 10.460000 1.600000 10.750000 1.645000 ;
      RECT 11.940000 0.735000 12.230000 0.780000 ;
      RECT 11.940000 0.920000 12.230000 0.965000 ;
  END
END sky130_fd_sc_hd__sedfxtp_4
MACRO sky130_fd_sc_hd__tap_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tap_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.265000 0.375000 0.810000 ;
      LAYER pwell ;
        RECT 0.145000 0.320000 0.315000 0.845000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.470000 0.375000 2.455000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
END sky130_fd_sc_hd__tap_1
MACRO sky130_fd_sc_hd__tap_2
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tap_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.920000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.920000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.265000 0.835000 0.810000 ;
      LAYER pwell ;
        RECT 0.145000 0.320000 0.775000 0.845000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.470000 0.835000 2.455000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 1.110000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.920000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.920000 0.085000 ;
      RECT 0.000000  2.635000 0.920000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
  END
END sky130_fd_sc_hd__tap_2
MACRO sky130_fd_sc_hd__tapvgnd2_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tapvgnd2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
      LAYER pwell ;
        RECT 0.145000 0.320000 0.315000 0.845000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.085000 1.755000 0.375000 1.985000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  1.470000 0.375000 2.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  1.785000 0.315000 1.955000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
END sky130_fd_sc_hd__tapvgnd2_1
MACRO sky130_fd_sc_hd__tapvgnd_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tapvgnd_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
      LAYER pwell ;
        RECT 0.145000 0.320000 0.315000 0.845000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.085000 2.095000 0.375000 2.325000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  1.470000 0.375000 2.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.125000 0.315000 2.295000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
END sky130_fd_sc_hd__tapvgnd_1
MACRO sky130_fd_sc_hd__tapvpwrvgnd_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tapvpwrvgnd_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
      LAYER pwell ;
        RECT 0.145000 0.320000 0.315000 0.845000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 2.910000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  1.470000 0.375000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
END sky130_fd_sc_hd__tapvpwrvgnd_1
MACRO sky130_fd_sc_hd__xnor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.930000 1.075000 1.625000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.670000 1.445000 ;
        RECT 0.425000 1.445000 1.965000 1.615000 ;
        RECT 1.795000 1.075000 2.395000 1.245000 ;
        RECT 1.795000 1.245000 1.965000 1.445000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.525000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.265000 2.125000 2.645000 2.295000 ;
        RECT 2.475000 1.755000 3.135000 1.955000 ;
        RECT 2.475000 1.955000 2.645000 2.125000 ;
        RECT 2.815000 0.345000 3.135000 0.825000 ;
        RECT 2.965000 0.825000 3.135000 1.755000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.280000 0.550000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.785000 ;
      RECT 0.085000  1.785000 2.305000 1.955000 ;
      RECT 0.085000  2.125000 0.385000 2.635000 ;
      RECT 0.555000  1.955000 0.885000 2.465000 ;
      RECT 1.055000  0.085000 1.225000 0.905000 ;
      RECT 1.055000  2.125000 1.685000 2.635000 ;
      RECT 1.395000  0.255000 1.725000 0.735000 ;
      RECT 1.395000  0.735000 2.645000 0.825000 ;
      RECT 1.395000  0.825000 2.305000 0.905000 ;
      RECT 1.895000  0.085000 2.245000 0.475000 ;
      RECT 2.135000  0.655000 2.645000 0.735000 ;
      RECT 2.135000  1.415000 2.795000 1.585000 ;
      RECT 2.135000  1.585000 2.305000 1.785000 ;
      RECT 2.415000  0.255000 2.645000 0.655000 ;
      RECT 2.625000  0.995000 2.795000 1.415000 ;
      RECT 2.815000  2.125000 3.115000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__xnor2_1
MACRO sky130_fd_sc_hd__xnor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.255000 1.075000 2.705000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.485000 1.075000 0.960000 1.285000 ;
        RECT 0.790000 1.285000 0.960000 1.445000 ;
        RECT 0.790000 1.445000 3.100000 1.615000 ;
        RECT 2.930000 1.075000 3.955000 1.285000 ;
        RECT 2.930000 1.285000 3.100000 1.445000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.913000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725000 1.795000 5.295000 1.965000 ;
        RECT 3.725000 1.965000 3.935000 2.125000 ;
        RECT 4.585000 0.305000 5.895000 0.475000 ;
        RECT 5.045000 1.415000 5.895000 1.625000 ;
        RECT 5.045000 1.625000 5.295000 1.795000 ;
        RECT 5.045000 1.965000 5.295000 2.125000 ;
        RECT 5.505000 0.475000 5.895000 1.415000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.645000 0.860000 0.895000 ;
      RECT 0.085000  0.895000 0.315000 1.785000 ;
      RECT 0.085000  1.785000 3.480000 1.955000 ;
      RECT 0.085000  1.955000 2.080000 1.965000 ;
      RECT 0.085000  1.965000 0.400000 2.465000 ;
      RECT 0.105000  0.255000 1.280000 0.475000 ;
      RECT 0.570000  2.135000 0.820000 2.635000 ;
      RECT 0.990000  1.965000 1.240000 2.465000 ;
      RECT 1.030000  0.475000 1.280000 0.725000 ;
      RECT 1.030000  0.725000 2.120000 0.905000 ;
      RECT 1.410000  2.135000 1.660000 2.635000 ;
      RECT 1.450000  0.085000 1.620000 0.555000 ;
      RECT 1.790000  0.255000 2.120000 0.725000 ;
      RECT 1.830000  1.965000 2.080000 2.465000 ;
      RECT 2.390000  2.125000 2.640000 2.465000 ;
      RECT 2.430000  0.085000 2.600000 0.905000 ;
      RECT 2.770000  0.255000 3.100000 0.725000 ;
      RECT 2.770000  0.725000 5.335000 0.905000 ;
      RECT 2.810000  2.135000 3.060000 2.635000 ;
      RECT 3.230000  2.125000 3.555000 2.295000 ;
      RECT 3.230000  2.295000 4.355000 2.465000 ;
      RECT 3.270000  0.085000 3.440000 0.555000 ;
      RECT 3.310000  1.455000 4.805000 1.625000 ;
      RECT 3.310000  1.625000 3.480000 1.785000 ;
      RECT 3.610000  0.255000 3.975000 0.725000 ;
      RECT 4.105000  2.135000 4.355000 2.295000 ;
      RECT 4.145000  0.085000 4.315000 0.555000 ;
      RECT 4.625000  2.135000 4.875000 2.635000 ;
      RECT 4.635000  1.075000 5.295000 1.245000 ;
      RECT 4.635000  1.245000 4.805000 1.455000 ;
      RECT 5.005000  0.645000 5.335000 0.725000 ;
      RECT 5.465000  1.795000 5.895000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.465000  2.125000 2.635000 2.295000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.385000  2.125000 3.555000 2.295000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 2.405000 2.095000 2.695000 2.140000 ;
      RECT 2.405000 2.140000 3.615000 2.280000 ;
      RECT 2.405000 2.280000 2.695000 2.325000 ;
      RECT 3.325000 2.095000 3.615000 2.140000 ;
      RECT 3.325000 2.280000 3.615000 2.325000 ;
  END
END sky130_fd_sc_hd__xnor2_2
MACRO sky130_fd_sc_hd__xnor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.175000 1.075000 5.390000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.490000 1.075000 1.855000 1.275000 ;
        RECT 1.685000 1.275000 1.855000 1.445000 ;
        RECT 1.685000 1.445000 5.730000 1.615000 ;
        RECT 5.560000 1.075000 7.430000 1.275000 ;
        RECT 5.560000 1.275000 5.730000 1.445000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.721000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.160000 1.785000  8.250000 2.045000 ;
        RECT 7.960000 1.445000 10.035000 1.665000 ;
        RECT 7.960000 1.665000  8.250000 1.785000 ;
        RECT 7.960000 2.045000  8.250000 2.465000 ;
        RECT 8.380000 0.645000 10.035000 0.905000 ;
        RECT 8.840000 1.665000  9.090000 2.465000 ;
        RECT 9.680000 1.665000 10.035000 2.465000 ;
        RECT 9.815000 0.905000 10.035000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.085000  0.645000  1.760000 0.905000 ;
      RECT 0.085000  0.905000  0.320000 1.445000 ;
      RECT 0.085000  1.445000  1.300000 1.615000 ;
      RECT 0.085000  1.615000  0.460000 2.465000 ;
      RECT 0.170000  0.255000  2.180000 0.475000 ;
      RECT 0.630000  1.835000  0.880000 2.635000 ;
      RECT 1.050000  1.615000  1.300000 1.785000 ;
      RECT 1.050000  1.785000  3.820000 2.005000 ;
      RECT 1.050000  2.005000  1.300000 2.465000 ;
      RECT 1.470000  2.175000  1.720000 2.635000 ;
      RECT 1.890000  2.005000  2.140000 2.465000 ;
      RECT 1.930000  0.475000  2.180000 0.725000 ;
      RECT 1.930000  0.725000  3.860000 0.905000 ;
      RECT 2.310000  2.175000  2.560000 2.635000 ;
      RECT 2.350000  0.085000  2.520000 0.555000 ;
      RECT 2.690000  0.255000  3.020000 0.725000 ;
      RECT 2.730000  2.005000  2.980000 2.465000 ;
      RECT 3.150000  2.175000  3.400000 2.635000 ;
      RECT 3.190000  0.085000  3.360000 0.555000 ;
      RECT 3.530000  0.255000  3.860000 0.725000 ;
      RECT 3.570000  2.005000  3.820000 2.465000 ;
      RECT 4.035000  0.085000  4.310000 0.905000 ;
      RECT 4.035000  1.785000  5.990000 2.005000 ;
      RECT 4.035000  2.005000  4.350000 2.465000 ;
      RECT 4.480000  0.255000  4.810000 0.725000 ;
      RECT 4.480000  0.725000  7.430000 0.735000 ;
      RECT 4.480000  0.735000  8.210000 0.905000 ;
      RECT 4.520000  2.175000  4.770000 2.635000 ;
      RECT 4.940000  2.005000  5.190000 2.465000 ;
      RECT 4.980000  0.085000  5.150000 0.555000 ;
      RECT 5.320000  0.255000  5.650000 0.725000 ;
      RECT 5.360000  2.175000  5.610000 2.635000 ;
      RECT 5.780000  2.005000  5.990000 2.215000 ;
      RECT 5.780000  2.215000  7.750000 2.465000 ;
      RECT 5.820000  0.085000  5.990000 0.555000 ;
      RECT 5.900000  1.445000  7.770000 1.615000 ;
      RECT 6.160000  0.255000  6.490000 0.725000 ;
      RECT 6.660000  0.085000  6.830000 0.555000 ;
      RECT 7.000000  0.255000  7.330000 0.725000 ;
      RECT 7.500000  0.085000  7.770000 0.555000 ;
      RECT 7.600000  1.075000  9.645000 1.275000 ;
      RECT 7.600000  1.275000  7.770000 1.445000 ;
      RECT 7.960000  0.305000  9.970000 0.475000 ;
      RECT 7.960000  0.475000  8.210000 0.735000 ;
      RECT 8.420000  1.835000  8.670000 2.635000 ;
      RECT 9.260000  1.835000  9.510000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  1.445000 1.235000 1.615000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  1.445000 6.295000 1.615000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
    LAYER met1 ;
      RECT 1.005000 1.415000 1.295000 1.460000 ;
      RECT 1.005000 1.460000 6.355000 1.600000 ;
      RECT 1.005000 1.600000 1.295000 1.645000 ;
      RECT 6.065000 1.415000 6.355000 1.460000 ;
      RECT 6.065000 1.600000 6.355000 1.645000 ;
  END
END sky130_fd_sc_hd__xnor2_4
MACRO sky130_fd_sc_hd__xnor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.045000 1.075000 7.455000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.225000 0.995000 6.395000 1.445000 ;
        RECT 6.225000 1.445000 6.805000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.615000 1.075000 2.180000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.345000 0.925000 ;
        RECT 0.085000 0.925000 0.330000 1.440000 ;
        RECT 0.085000 1.440000 0.365000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.500000  0.995000 0.705000 1.325000 ;
      RECT 0.515000  0.085000 0.765000 0.525000 ;
      RECT 0.530000  0.695000 1.105000 0.865000 ;
      RECT 0.530000  0.865000 0.705000 0.995000 ;
      RECT 0.535000  1.325000 0.705000 1.875000 ;
      RECT 0.535000  1.875000 1.220000 2.045000 ;
      RECT 0.535000  2.215000 0.870000 2.635000 ;
      RECT 0.935000  0.255000 2.505000 0.425000 ;
      RECT 0.935000  0.425000 1.105000 0.695000 ;
      RECT 0.935000  1.535000 2.520000 1.705000 ;
      RECT 1.050000  2.045000 1.220000 2.235000 ;
      RECT 1.050000  2.235000 2.520000 2.405000 ;
      RECT 1.275000  0.595000 1.445000 1.535000 ;
      RECT 1.560000  1.895000 4.060000 2.065000 ;
      RECT 1.745000  0.625000 2.965000 0.795000 ;
      RECT 1.745000  0.795000 2.125000 0.905000 ;
      RECT 2.070000  0.425000 2.505000 0.455000 ;
      RECT 2.350000  0.995000 2.625000 1.325000 ;
      RECT 2.350000  1.325000 2.520000 1.535000 ;
      RECT 2.675000  0.285000 3.305000 0.455000 ;
      RECT 2.690000  1.525000 3.075000 1.695000 ;
      RECT 2.795000  0.795000 2.965000 1.375000 ;
      RECT 2.795000  1.375000 3.075000 1.525000 ;
      RECT 3.135000  0.455000 3.305000 1.035000 ;
      RECT 3.135000  1.035000 3.415000 1.205000 ;
      RECT 3.225000  2.235000 3.555000 2.635000 ;
      RECT 3.245000  1.205000 3.415000 1.895000 ;
      RECT 3.475000  0.085000 3.645000 0.865000 ;
      RECT 3.645000  1.445000 4.065000 1.715000 ;
      RECT 3.825000  0.415000 4.065000 1.445000 ;
      RECT 3.890000  2.065000 4.060000 2.275000 ;
      RECT 3.890000  2.275000 6.985000 2.445000 ;
      RECT 4.245000  0.265000 4.655000 0.485000 ;
      RECT 4.245000  0.485000 4.455000 0.595000 ;
      RECT 4.245000  0.595000 4.415000 2.105000 ;
      RECT 4.585000  0.720000 4.995000 0.825000 ;
      RECT 4.585000  0.825000 4.795000 0.890000 ;
      RECT 4.585000  0.890000 4.755000 2.275000 ;
      RECT 4.625000  0.655000 4.995000 0.720000 ;
      RECT 4.825000  0.320000 4.995000 0.655000 ;
      RECT 4.935000  1.445000 5.715000 1.615000 ;
      RECT 4.935000  1.615000 5.350000 2.045000 ;
      RECT 4.950000  0.995000 5.375000 1.270000 ;
      RECT 5.165000  0.630000 5.375000 0.995000 ;
      RECT 5.545000  0.255000 6.690000 0.425000 ;
      RECT 5.545000  0.425000 5.715000 1.445000 ;
      RECT 5.885000  0.595000 6.055000 1.935000 ;
      RECT 5.885000  1.935000 8.195000 2.105000 ;
      RECT 6.225000  0.425000 6.690000 0.465000 ;
      RECT 6.565000  0.730000 6.770000 0.945000 ;
      RECT 6.565000  0.945000 6.875000 1.275000 ;
      RECT 6.975000  1.495000 7.795000 1.705000 ;
      RECT 7.015000  0.295000 7.305000 0.735000 ;
      RECT 7.015000  0.735000 7.795000 0.750000 ;
      RECT 7.055000  0.750000 7.795000 0.905000 ;
      RECT 7.395000  2.275000 7.730000 2.635000 ;
      RECT 7.475000  0.085000 7.645000 0.565000 ;
      RECT 7.625000  0.905000 7.795000 0.995000 ;
      RECT 7.625000  0.995000 7.855000 1.325000 ;
      RECT 7.625000  1.325000 7.795000 1.495000 ;
      RECT 7.710000  1.875000 8.195000 1.935000 ;
      RECT 7.895000  0.255000 8.195000 0.585000 ;
      RECT 7.900000  2.105000 8.195000 2.465000 ;
      RECT 8.025000  0.585000 8.195000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  1.445000 3.075000 1.615000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  0.765000 3.995000 0.935000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  0.425000 4.455000 0.595000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  0.765000 5.375000 0.935000 ;
      RECT 5.205000  1.445000 5.375000 1.615000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  0.765000 6.755000 0.935000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  0.425000 7.215000 0.595000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
    LAYER met1 ;
      RECT 2.845000 1.415000 3.135000 1.460000 ;
      RECT 2.845000 1.460000 5.435000 1.600000 ;
      RECT 2.845000 1.600000 3.135000 1.645000 ;
      RECT 3.765000 0.735000 4.055000 0.780000 ;
      RECT 3.765000 0.780000 6.815000 0.920000 ;
      RECT 3.765000 0.920000 4.055000 0.965000 ;
      RECT 4.225000 0.395000 4.515000 0.440000 ;
      RECT 4.225000 0.440000 7.275000 0.580000 ;
      RECT 4.225000 0.580000 4.515000 0.625000 ;
      RECT 5.145000 0.735000 5.435000 0.780000 ;
      RECT 5.145000 0.920000 5.435000 0.965000 ;
      RECT 5.145000 1.415000 5.435000 1.460000 ;
      RECT 5.145000 1.600000 5.435000 1.645000 ;
      RECT 6.525000 0.735000 6.815000 0.780000 ;
      RECT 6.525000 0.920000 6.815000 0.965000 ;
      RECT 6.985000 0.395000 7.275000 0.440000 ;
      RECT 6.985000 0.580000 7.275000 0.625000 ;
  END
END sky130_fd_sc_hd__xnor3_1
MACRO sky130_fd_sc_hd__xnor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.505000 1.075000 7.915000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.685000 0.995000 6.855000 1.445000 ;
        RECT 6.685000 1.445000 7.265000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.075000 2.640000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.350000 0.805000 0.925000 ;
        RECT 0.545000 0.925000 0.790000 1.440000 ;
        RECT 0.545000 1.440000 0.825000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.930000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.085000  0.085000 0.375000 0.735000 ;
      RECT 0.085000  1.490000 0.375000 2.635000 ;
      RECT 0.960000  0.995000 1.165000 1.325000 ;
      RECT 0.975000  0.085000 1.225000 0.525000 ;
      RECT 0.990000  0.695000 1.565000 0.865000 ;
      RECT 0.990000  0.865000 1.165000 0.995000 ;
      RECT 0.995000  1.325000 1.165000 1.875000 ;
      RECT 0.995000  1.875000 1.680000 2.045000 ;
      RECT 0.995000  2.215000 1.330000 2.635000 ;
      RECT 1.395000  0.255000 2.965000 0.425000 ;
      RECT 1.395000  0.425000 1.565000 0.695000 ;
      RECT 1.395000  1.535000 2.980000 1.705000 ;
      RECT 1.510000  2.045000 1.680000 2.235000 ;
      RECT 1.510000  2.235000 2.980000 2.405000 ;
      RECT 1.735000  0.595000 1.905000 1.535000 ;
      RECT 2.020000  1.895000 4.520000 2.065000 ;
      RECT 2.205000  0.625000 3.425000 0.795000 ;
      RECT 2.205000  0.795000 2.585000 0.905000 ;
      RECT 2.530000  0.425000 2.965000 0.455000 ;
      RECT 2.810000  0.995000 3.085000 1.325000 ;
      RECT 2.810000  1.325000 2.980000 1.535000 ;
      RECT 3.135000  0.285000 3.765000 0.455000 ;
      RECT 3.150000  1.525000 3.535000 1.695000 ;
      RECT 3.255000  0.795000 3.425000 1.375000 ;
      RECT 3.255000  1.375000 3.535000 1.525000 ;
      RECT 3.595000  0.455000 3.765000 1.035000 ;
      RECT 3.595000  1.035000 3.875000 1.205000 ;
      RECT 3.685000  2.235000 4.015000 2.635000 ;
      RECT 3.705000  1.205000 3.875000 1.895000 ;
      RECT 3.935000  0.085000 4.105000 0.865000 ;
      RECT 4.105000  1.445000 4.525000 1.715000 ;
      RECT 4.285000  0.415000 4.525000 1.445000 ;
      RECT 4.350000  2.065000 4.520000 2.275000 ;
      RECT 4.350000  2.275000 7.445000 2.445000 ;
      RECT 4.705000  0.265000 5.115000 0.485000 ;
      RECT 4.705000  0.485000 4.915000 0.595000 ;
      RECT 4.705000  0.595000 4.875000 2.105000 ;
      RECT 5.045000  0.720000 5.455000 0.825000 ;
      RECT 5.045000  0.825000 5.255000 0.890000 ;
      RECT 5.045000  0.890000 5.215000 2.275000 ;
      RECT 5.085000  0.655000 5.455000 0.720000 ;
      RECT 5.285000  0.320000 5.455000 0.655000 ;
      RECT 5.395000  1.445000 6.175000 1.615000 ;
      RECT 5.395000  1.615000 5.810000 2.045000 ;
      RECT 5.410000  0.995000 5.835000 1.270000 ;
      RECT 5.625000  0.630000 5.835000 0.995000 ;
      RECT 6.005000  0.255000 7.150000 0.425000 ;
      RECT 6.005000  0.425000 6.175000 1.445000 ;
      RECT 6.345000  0.595000 6.515000 1.935000 ;
      RECT 6.345000  1.935000 8.655000 2.105000 ;
      RECT 6.685000  0.425000 7.150000 0.465000 ;
      RECT 7.025000  0.730000 7.230000 0.945000 ;
      RECT 7.025000  0.945000 7.335000 1.275000 ;
      RECT 7.435000  1.495000 8.255000 1.705000 ;
      RECT 7.475000  0.295000 7.765000 0.735000 ;
      RECT 7.475000  0.735000 8.255000 0.750000 ;
      RECT 7.515000  0.750000 8.255000 0.905000 ;
      RECT 7.855000  2.275000 8.190000 2.635000 ;
      RECT 7.935000  0.085000 8.105000 0.565000 ;
      RECT 8.085000  0.905000 8.255000 0.995000 ;
      RECT 8.085000  0.995000 8.315000 1.325000 ;
      RECT 8.085000  1.325000 8.255000 1.495000 ;
      RECT 8.170000  1.875000 8.655000 1.935000 ;
      RECT 8.355000  0.255000 8.655000 0.585000 ;
      RECT 8.360000  2.105000 8.655000 2.465000 ;
      RECT 8.485000  0.585000 8.655000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  1.445000 3.535000 1.615000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  0.765000 4.455000 0.935000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  0.425000 4.915000 0.595000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  0.765000 5.835000 0.935000 ;
      RECT 5.665000  1.445000 5.835000 1.615000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  0.765000 7.215000 0.935000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  0.425000 7.675000 0.595000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
    LAYER met1 ;
      RECT 3.305000 1.415000 3.595000 1.460000 ;
      RECT 3.305000 1.460000 5.895000 1.600000 ;
      RECT 3.305000 1.600000 3.595000 1.645000 ;
      RECT 4.225000 0.735000 4.515000 0.780000 ;
      RECT 4.225000 0.780000 7.275000 0.920000 ;
      RECT 4.225000 0.920000 4.515000 0.965000 ;
      RECT 4.685000 0.395000 4.975000 0.440000 ;
      RECT 4.685000 0.440000 7.735000 0.580000 ;
      RECT 4.685000 0.580000 4.975000 0.625000 ;
      RECT 5.605000 0.735000 5.895000 0.780000 ;
      RECT 5.605000 0.920000 5.895000 0.965000 ;
      RECT 5.605000 1.415000 5.895000 1.460000 ;
      RECT 5.605000 1.600000 5.895000 1.645000 ;
      RECT 6.985000 0.735000 7.275000 0.780000 ;
      RECT 6.985000 0.920000 7.275000 0.965000 ;
      RECT 7.445000 0.395000 7.735000 0.440000 ;
      RECT 7.445000 0.580000 7.735000 0.625000 ;
  END
END sky130_fd_sc_hd__xnor3_2
MACRO sky130_fd_sc_hd__xnor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.425000 1.075000 8.835000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.605000 0.995000 7.775000 1.445000 ;
        RECT 7.605000 1.445000 8.185000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.995000 1.075000 3.560000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 0.375000 0.875000 0.995000 ;
        RECT 0.625000 0.995000 1.710000 1.325000 ;
        RECT 0.625000 1.325000 0.955000 2.425000 ;
        RECT 1.465000 0.350000 1.725000 0.925000 ;
        RECT 1.465000 0.925000 1.710000 0.995000 ;
        RECT 1.465000 1.325000 1.710000 1.440000 ;
        RECT 1.465000 1.440000 1.745000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.285000  0.085000 0.455000 0.735000 ;
      RECT 0.285000  1.490000 0.455000 2.635000 ;
      RECT 1.125000  0.085000 1.295000 0.735000 ;
      RECT 1.125000  1.495000 1.295000 2.635000 ;
      RECT 1.880000  0.995000 2.085000 1.325000 ;
      RECT 1.895000  0.085000 2.145000 0.525000 ;
      RECT 1.910000  0.695000 2.485000 0.865000 ;
      RECT 1.910000  0.865000 2.085000 0.995000 ;
      RECT 1.915000  1.325000 2.085000 1.875000 ;
      RECT 1.915000  1.875000 2.600000 2.045000 ;
      RECT 1.915000  2.215000 2.250000 2.635000 ;
      RECT 2.315000  0.255000 3.885000 0.425000 ;
      RECT 2.315000  0.425000 2.485000 0.695000 ;
      RECT 2.315000  1.535000 3.900000 1.705000 ;
      RECT 2.430000  2.045000 2.600000 2.235000 ;
      RECT 2.430000  2.235000 3.900000 2.405000 ;
      RECT 2.655000  0.595000 2.825000 1.535000 ;
      RECT 2.940000  1.895000 5.440000 2.065000 ;
      RECT 3.125000  0.625000 4.345000 0.795000 ;
      RECT 3.125000  0.795000 3.505000 0.905000 ;
      RECT 3.450000  0.425000 3.885000 0.455000 ;
      RECT 3.730000  0.995000 4.005000 1.325000 ;
      RECT 3.730000  1.325000 3.900000 1.535000 ;
      RECT 4.055000  0.285000 4.685000 0.455000 ;
      RECT 4.070000  1.525000 4.455000 1.695000 ;
      RECT 4.175000  0.795000 4.345000 1.375000 ;
      RECT 4.175000  1.375000 4.455000 1.525000 ;
      RECT 4.515000  0.455000 4.685000 1.035000 ;
      RECT 4.515000  1.035000 4.795000 1.205000 ;
      RECT 4.605000  2.235000 4.935000 2.635000 ;
      RECT 4.625000  1.205000 4.795000 1.895000 ;
      RECT 4.855000  0.085000 5.025000 0.865000 ;
      RECT 5.025000  1.445000 5.445000 1.715000 ;
      RECT 5.205000  0.415000 5.445000 1.445000 ;
      RECT 5.270000  2.065000 5.440000 2.275000 ;
      RECT 5.270000  2.275000 8.365000 2.445000 ;
      RECT 5.625000  0.265000 6.035000 0.485000 ;
      RECT 5.625000  0.485000 5.835000 0.595000 ;
      RECT 5.625000  0.595000 5.795000 2.105000 ;
      RECT 5.965000  0.720000 6.375000 0.825000 ;
      RECT 5.965000  0.825000 6.175000 0.890000 ;
      RECT 5.965000  0.890000 6.135000 2.275000 ;
      RECT 6.005000  0.655000 6.375000 0.720000 ;
      RECT 6.205000  0.320000 6.375000 0.655000 ;
      RECT 6.315000  1.445000 7.095000 1.615000 ;
      RECT 6.315000  1.615000 6.730000 2.045000 ;
      RECT 6.330000  0.995000 6.755000 1.270000 ;
      RECT 6.545000  0.630000 6.755000 0.995000 ;
      RECT 6.925000  0.255000 8.070000 0.425000 ;
      RECT 6.925000  0.425000 7.095000 1.445000 ;
      RECT 7.265000  0.595000 7.435000 1.935000 ;
      RECT 7.265000  1.935000 9.575000 2.105000 ;
      RECT 7.605000  0.425000 8.070000 0.465000 ;
      RECT 7.945000  0.730000 8.150000 0.945000 ;
      RECT 7.945000  0.945000 8.255000 1.275000 ;
      RECT 8.355000  1.495000 9.175000 1.705000 ;
      RECT 8.395000  0.295000 8.685000 0.735000 ;
      RECT 8.395000  0.735000 9.175000 0.750000 ;
      RECT 8.435000  0.750000 9.175000 0.905000 ;
      RECT 8.775000  2.275000 9.110000 2.635000 ;
      RECT 8.855000  0.085000 9.025000 0.565000 ;
      RECT 9.005000  0.905000 9.175000 0.995000 ;
      RECT 9.005000  0.995000 9.235000 1.325000 ;
      RECT 9.005000  1.325000 9.175000 1.495000 ;
      RECT 9.090000  1.875000 9.575000 1.935000 ;
      RECT 9.275000  0.255000 9.575000 0.585000 ;
      RECT 9.280000  2.105000 9.575000 2.465000 ;
      RECT 9.405000  0.585000 9.575000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  1.445000 4.455000 1.615000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  0.765000 5.375000 0.935000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  0.425000 5.835000 0.595000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  0.765000 6.755000 0.935000 ;
      RECT 6.585000  1.445000 6.755000 1.615000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  0.765000 8.135000 0.935000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  0.425000 8.595000 0.595000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 4.225000 1.415000 4.515000 1.460000 ;
      RECT 4.225000 1.460000 6.815000 1.600000 ;
      RECT 4.225000 1.600000 4.515000 1.645000 ;
      RECT 5.145000 0.735000 5.435000 0.780000 ;
      RECT 5.145000 0.780000 8.195000 0.920000 ;
      RECT 5.145000 0.920000 5.435000 0.965000 ;
      RECT 5.605000 0.395000 5.895000 0.440000 ;
      RECT 5.605000 0.440000 8.655000 0.580000 ;
      RECT 5.605000 0.580000 5.895000 0.625000 ;
      RECT 6.525000 0.735000 6.815000 0.780000 ;
      RECT 6.525000 0.920000 6.815000 0.965000 ;
      RECT 6.525000 1.415000 6.815000 1.460000 ;
      RECT 6.525000 1.600000 6.815000 1.645000 ;
      RECT 7.905000 0.735000 8.195000 0.780000 ;
      RECT 7.905000 0.920000 8.195000 0.965000 ;
      RECT 8.365000 0.395000 8.655000 0.440000 ;
      RECT 8.365000 0.580000 8.655000 0.625000 ;
  END
END sky130_fd_sc_hd__xnor3_4
MACRO sky130_fd_sc_hd__xor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.840000 1.075000 1.390000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.670000 1.445000 ;
        RECT 0.425000 1.445000 1.730000 1.615000 ;
        RECT 1.560000 1.075000 1.935000 1.245000 ;
        RECT 1.560000 1.245000 1.730000 1.445000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.800500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.720000 0.315000 2.675000 0.485000 ;
        RECT 2.505000 0.485000 2.675000 1.365000 ;
        RECT 2.505000 1.365000 3.135000 1.535000 ;
        RECT 2.815000 1.535000 3.135000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.655000 2.335000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.785000 ;
      RECT 0.085000  1.785000 0.465000 2.465000 ;
      RECT 0.135000  0.085000 0.465000 0.475000 ;
      RECT 0.635000  0.335000 0.805000 0.655000 ;
      RECT 0.975000  0.085000 1.305000 0.475000 ;
      RECT 1.055000  1.785000 1.225000 2.635000 ;
      RECT 1.395000  1.785000 2.635000 1.955000 ;
      RECT 1.395000  1.955000 1.725000 2.465000 ;
      RECT 1.895000  2.125000 2.065000 2.635000 ;
      RECT 2.105000  0.825000 2.335000 1.325000 ;
      RECT 2.235000  1.955000 2.635000 2.465000 ;
      RECT 2.845000  0.085000 3.135000 0.920000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__xor2_1
MACRO sky130_fd_sc_hd__xor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.075000 0.875000 1.275000 ;
        RECT 0.705000 1.275000 0.875000 1.445000 ;
        RECT 0.705000 1.445000 1.880000 1.615000 ;
        RECT 1.710000 1.075000 3.230000 1.275000 ;
        RECT 1.710000 1.275000 1.880000 1.445000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.075000 1.540000 1.275000 ;
      LAYER mcon ;
        RECT 1.065000 1.105000 1.235000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.420000 1.075000 4.090000 1.275000 ;
      LAYER mcon ;
        RECT 3.825000 1.105000 3.995000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.005000 1.075000 1.295000 1.120000 ;
        RECT 1.005000 1.120000 4.055000 1.260000 ;
        RECT 1.005000 1.260000 1.295000 1.305000 ;
        RECT 3.765000 1.075000 4.055000 1.120000 ;
        RECT 3.765000 1.260000 4.055000 1.305000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.656750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.625000 0.645000 3.955000 0.725000 ;
        RECT 3.625000 0.725000 5.895000 0.905000 ;
        RECT 4.985000 0.645000 5.315000 0.725000 ;
        RECT 5.025000 1.415000 5.895000 1.625000 ;
        RECT 5.025000 1.625000 5.275000 2.125000 ;
        RECT 5.485000 0.905000 5.895000 1.415000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.120000  0.725000 1.700000 0.905000 ;
      RECT 0.120000  0.905000 0.290000 1.785000 ;
      RECT 0.120000  1.785000 2.220000 1.955000 ;
      RECT 0.120000  2.135000 0.400000 2.465000 ;
      RECT 0.145000  2.125000 0.315000 2.135000 ;
      RECT 0.190000  0.085000 0.360000 0.555000 ;
      RECT 0.530000  0.255000 0.860000 0.725000 ;
      RECT 0.570000  2.135000 0.820000 2.635000 ;
      RECT 0.990000  2.135000 1.240000 2.295000 ;
      RECT 0.990000  2.295000 2.080000 2.465000 ;
      RECT 1.030000  0.085000 1.200000 0.555000 ;
      RECT 1.065000  2.125000 1.235000 2.135000 ;
      RECT 1.370000  0.255000 1.700000 0.725000 ;
      RECT 1.410000  1.955000 1.660000 2.125000 ;
      RECT 1.830000  2.135000 2.080000 2.295000 ;
      RECT 1.870000  0.085000 2.040000 0.555000 ;
      RECT 2.050000  1.445000 4.785000 1.615000 ;
      RECT 2.050000  1.615000 2.220000 1.785000 ;
      RECT 2.285000  2.125000 2.600000 2.465000 ;
      RECT 2.310000  0.255000 2.640000 0.725000 ;
      RECT 2.310000  0.725000 3.400000 0.905000 ;
      RECT 2.390000  1.785000 4.855000 1.955000 ;
      RECT 2.390000  1.955000 2.600000 2.125000 ;
      RECT 2.770000  2.135000 3.020000 2.635000 ;
      RECT 2.810000  0.085000 2.980000 0.555000 ;
      RECT 3.150000  0.255000 4.380000 0.475000 ;
      RECT 3.150000  0.475000 3.400000 0.725000 ;
      RECT 3.190000  1.955000 3.440000 2.465000 ;
      RECT 3.610000  2.135000 3.915000 2.635000 ;
      RECT 4.085000  1.955000 4.855000 2.295000 ;
      RECT 4.085000  2.295000 5.695000 2.465000 ;
      RECT 4.615000  1.075000 5.275000 1.245000 ;
      RECT 4.615000  1.245000 4.785000 1.445000 ;
      RECT 4.645000  0.085000 4.815000 0.555000 ;
      RECT 5.445000  1.795000 5.695000 2.295000 ;
      RECT 5.485000  0.085000 5.655000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 0.085000 2.095000 0.375000 2.140000 ;
      RECT 0.085000 2.140000 1.295000 2.280000 ;
      RECT 0.085000 2.280000 0.375000 2.325000 ;
      RECT 1.005000 2.095000 1.295000 2.140000 ;
      RECT 1.005000 2.280000 1.295000 2.325000 ;
  END
END sky130_fd_sc_hd__xor2_2
MACRO sky130_fd_sc_hd__xor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 2.800000 1.275000 ;
        RECT 2.630000 1.275000 2.800000 1.445000 ;
        RECT 2.630000 1.445000 6.165000 1.615000 ;
        RECT 5.995000 1.075000 7.370000 1.275000 ;
        RECT 5.995000 1.275000 6.165000 1.445000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.075000 5.000000 1.105000 ;
        RECT 2.970000 1.105000 5.740000 1.275000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.524450 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165000 0.645000 5.580000 0.905000 ;
        RECT 5.150000 0.905000 5.580000 0.935000 ;
      LAYER mcon ;
        RECT 5.205000 0.765000 5.375000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.850000 0.725000  8.630000 0.735000 ;
        RECT 7.850000 0.735000 10.035000 0.905000 ;
        RECT 7.850000 0.905000  8.305000 0.935000 ;
        RECT 7.880000 1.445000 10.035000 1.625000 ;
        RECT 7.880000 1.625000  9.010000 1.665000 ;
        RECT 7.880000 1.665000  8.170000 2.125000 ;
        RECT 8.300000 0.255000  8.630000 0.725000 ;
        RECT 8.760000 1.665000  9.010000 2.125000 ;
        RECT 9.140000 0.255000  9.470000 0.735000 ;
        RECT 9.600000 1.625000 10.035000 2.465000 ;
        RECT 9.735000 0.905000 10.035000 1.445000 ;
      LAYER mcon ;
        RECT 7.965000 0.765000 8.135000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.145000 0.735000 5.435000 0.780000 ;
        RECT 5.145000 0.780000 8.195000 0.920000 ;
        RECT 5.145000 0.920000 5.435000 0.965000 ;
        RECT 7.905000 0.735000 8.195000 0.780000 ;
        RECT 7.905000 0.920000 8.195000 0.965000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.085000  0.085000  0.360000 0.565000 ;
      RECT 0.085000  0.735000  3.380000 0.905000 ;
      RECT 0.085000  0.905000  0.255000 1.445000 ;
      RECT 0.085000  1.445000  2.420000 1.615000 ;
      RECT 0.085000  1.785000  2.080000 2.005000 ;
      RECT 0.085000  2.005000  0.400000 2.465000 ;
      RECT 0.530000  0.255000  0.860000 0.725000 ;
      RECT 0.530000  0.725000  3.380000 0.735000 ;
      RECT 0.570000  2.175000  0.820000 2.635000 ;
      RECT 0.990000  2.005000  1.240000 2.465000 ;
      RECT 1.030000  0.085000  1.200000 0.555000 ;
      RECT 1.370000  0.255000  1.700000 0.725000 ;
      RECT 1.410000  2.175000  1.660000 2.635000 ;
      RECT 1.830000  2.005000  2.080000 2.295000 ;
      RECT 1.830000  2.295000  3.760000 2.465000 ;
      RECT 1.870000  0.085000  2.040000 0.555000 ;
      RECT 2.210000  0.255000  2.540000 0.725000 ;
      RECT 2.250000  1.615000  2.420000 1.785000 ;
      RECT 2.250000  1.785000  3.340000 1.955000 ;
      RECT 2.250000  1.955000  2.500000 2.125000 ;
      RECT 2.670000  2.125000  2.920000 2.295000 ;
      RECT 2.710000  0.085000  2.880000 0.555000 ;
      RECT 3.050000  0.255000  3.380000 0.725000 ;
      RECT 3.090000  1.955000  3.340000 2.125000 ;
      RECT 3.510000  1.795000  3.760000 2.295000 ;
      RECT 3.550000  0.085000  3.820000 0.895000 ;
      RECT 3.990000  0.255000  6.000000 0.475000 ;
      RECT 4.030000  1.785000  7.640000 2.005000 ;
      RECT 4.030000  2.005000  4.280000 2.465000 ;
      RECT 4.450000  2.175000  4.700000 2.635000 ;
      RECT 4.870000  2.005000  5.120000 2.465000 ;
      RECT 5.290000  2.175000  5.540000 2.635000 ;
      RECT 5.710000  2.005000  5.960000 2.465000 ;
      RECT 5.750000  0.475000  6.000000 0.725000 ;
      RECT 5.750000  0.725000  7.680000 0.905000 ;
      RECT 6.130000  2.175000  6.380000 2.635000 ;
      RECT 6.170000  0.085000  6.340000 0.555000 ;
      RECT 6.510000  0.255000  6.840000 0.725000 ;
      RECT 6.550000  1.455000  6.800000 1.785000 ;
      RECT 6.550000  2.005000  6.800000 2.465000 ;
      RECT 6.970000  2.175000  7.220000 2.635000 ;
      RECT 7.010000  0.085000  7.180000 0.555000 ;
      RECT 7.260000  1.445000  7.710000 1.615000 ;
      RECT 7.350000  0.255000  7.680000 0.725000 ;
      RECT 7.390000  2.005000  7.640000 2.295000 ;
      RECT 7.390000  2.295000  9.430000 2.465000 ;
      RECT 7.540000  1.105000  9.565000 1.275000 ;
      RECT 7.540000  1.275000  7.710000 1.445000 ;
      RECT 7.960000  0.085000  8.130000 0.555000 ;
      RECT 8.340000  1.835000  8.590000 2.295000 ;
      RECT 8.540000  1.075000  9.565000 1.105000 ;
      RECT 8.800000  0.085000  8.970000 0.555000 ;
      RECT 9.180000  1.795000  9.430000 2.295000 ;
      RECT 9.640000  0.085000  9.810000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  1.445000 2.155000 1.615000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  1.445000 7.675000 1.615000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
    LAYER met1 ;
      RECT 1.925000 1.415000 2.215000 1.460000 ;
      RECT 1.925000 1.460000 7.735000 1.600000 ;
      RECT 1.925000 1.600000 2.215000 1.645000 ;
      RECT 7.445000 1.415000 7.735000 1.460000 ;
      RECT 7.445000 1.600000 7.735000 1.645000 ;
  END
END sky130_fd_sc_hd__xor2_4
MACRO sky130_fd_sc_hd__xor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.505000 1.075000 7.915000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.685000 0.995000 6.855000 1.445000 ;
        RECT 6.685000 1.445000 7.265000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.860000 0.995000 2.495000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.590000 0.925000 ;
        RECT 0.085000 0.925000 0.400000 1.440000 ;
        RECT 0.085000 1.440000 0.610000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.930000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.750000  0.995000 0.950000 1.325000 ;
      RECT 0.760000  0.085000 1.010000 0.525000 ;
      RECT 0.780000  0.695000 1.350000 0.865000 ;
      RECT 0.780000  0.865000 0.950000 0.995000 ;
      RECT 0.780000  1.325000 0.950000 1.875000 ;
      RECT 0.780000  1.875000 1.470000 2.045000 ;
      RECT 0.780000  2.215000 1.115000 2.635000 ;
      RECT 1.180000  0.255000 2.740000 0.425000 ;
      RECT 1.180000  0.425000 1.350000 0.695000 ;
      RECT 1.185000  1.535000 2.835000 1.705000 ;
      RECT 1.300000  2.045000 1.470000 2.235000 ;
      RECT 1.300000  2.235000 2.895000 2.405000 ;
      RECT 1.520000  0.595000 1.690000 1.535000 ;
      RECT 1.870000  1.895000 3.175000 2.065000 ;
      RECT 1.970000  0.655000 3.080000 0.825000 ;
      RECT 2.390000  0.425000 2.740000 0.455000 ;
      RECT 2.665000  0.995000 2.940000 1.325000 ;
      RECT 2.665000  1.325000 2.835000 1.535000 ;
      RECT 2.910000  0.255000 3.760000 0.425000 ;
      RECT 2.910000  0.425000 3.080000 0.655000 ;
      RECT 3.005000  1.525000 3.535000 1.695000 ;
      RECT 3.005000  1.695000 3.175000 1.895000 ;
      RECT 3.110000  2.235000 3.515000 2.405000 ;
      RECT 3.250000  0.595000 3.420000 1.375000 ;
      RECT 3.250000  1.375000 3.535000 1.525000 ;
      RECT 3.345000  1.895000 4.520000 2.065000 ;
      RECT 3.345000  2.065000 3.515000 2.235000 ;
      RECT 3.590000  0.425000 3.760000 1.035000 ;
      RECT 3.590000  1.035000 3.875000 1.205000 ;
      RECT 3.685000  2.235000 4.015000 2.635000 ;
      RECT 3.705000  1.205000 3.875000 1.895000 ;
      RECT 3.930000  0.085000 4.100000 0.865000 ;
      RECT 4.105000  1.445000 4.520000 1.715000 ;
      RECT 4.280000  0.415000 4.520000 1.445000 ;
      RECT 4.350000  2.065000 4.520000 2.275000 ;
      RECT 4.350000  2.275000 7.445000 2.445000 ;
      RECT 4.695000  0.265000 5.110000 0.485000 ;
      RECT 4.695000  0.485000 4.915000 0.595000 ;
      RECT 4.695000  0.595000 4.865000 2.105000 ;
      RECT 5.035000  0.720000 5.450000 0.825000 ;
      RECT 5.035000  0.825000 5.255000 0.890000 ;
      RECT 5.035000  0.890000 5.205000 2.275000 ;
      RECT 5.085000  0.655000 5.450000 0.720000 ;
      RECT 5.280000  0.320000 5.450000 0.655000 ;
      RECT 5.395000  1.445000 6.175000 1.615000 ;
      RECT 5.395000  1.615000 5.810000 2.045000 ;
      RECT 5.410000  0.995000 5.835000 1.270000 ;
      RECT 5.620000  0.630000 5.835000 0.995000 ;
      RECT 6.005000  0.255000 7.150000 0.425000 ;
      RECT 6.005000  0.425000 6.175000 1.445000 ;
      RECT 6.345000  0.595000 6.515000 1.935000 ;
      RECT 6.345000  1.935000 8.655000 2.105000 ;
      RECT 6.685000  0.425000 7.150000 0.465000 ;
      RECT 7.025000  0.730000 7.230000 0.945000 ;
      RECT 7.025000  0.945000 7.335000 1.275000 ;
      RECT 7.435000  1.495000 8.255000 1.705000 ;
      RECT 7.475000  0.295000 7.765000 0.735000 ;
      RECT 7.475000  0.735000 8.255000 0.750000 ;
      RECT 7.515000  0.750000 8.255000 0.905000 ;
      RECT 7.855000  2.275000 8.190000 2.635000 ;
      RECT 7.935000  0.085000 8.105000 0.565000 ;
      RECT 8.085000  0.905000 8.255000 0.995000 ;
      RECT 8.085000  0.995000 8.315000 1.325000 ;
      RECT 8.085000  1.325000 8.255000 1.495000 ;
      RECT 8.170000  1.875000 8.655000 1.935000 ;
      RECT 8.355000  0.255000 8.655000 0.585000 ;
      RECT 8.360000  2.105000 8.655000 2.465000 ;
      RECT 8.485000  0.585000 8.655000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  1.445000 3.535000 1.615000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  0.765000 4.455000 0.935000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  0.425000 4.915000 0.595000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  0.765000 5.835000 0.935000 ;
      RECT 5.665000  1.445000 5.835000 1.615000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  0.765000 7.215000 0.935000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  0.425000 7.675000 0.595000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
    LAYER met1 ;
      RECT 3.305000 1.415000 3.595000 1.460000 ;
      RECT 3.305000 1.460000 5.895000 1.600000 ;
      RECT 3.305000 1.600000 3.595000 1.645000 ;
      RECT 4.225000 0.735000 4.515000 0.780000 ;
      RECT 4.225000 0.780000 7.275000 0.920000 ;
      RECT 4.225000 0.920000 4.515000 0.965000 ;
      RECT 4.685000 0.395000 4.975000 0.440000 ;
      RECT 4.685000 0.440000 7.735000 0.580000 ;
      RECT 4.685000 0.580000 4.975000 0.625000 ;
      RECT 5.605000 0.735000 5.895000 0.780000 ;
      RECT 5.605000 0.920000 5.895000 0.965000 ;
      RECT 5.605000 1.415000 5.895000 1.460000 ;
      RECT 5.605000 1.600000 5.895000 1.645000 ;
      RECT 6.985000 0.735000 7.275000 0.780000 ;
      RECT 6.985000 0.920000 7.275000 0.965000 ;
      RECT 7.445000 0.395000 7.735000 0.440000 ;
      RECT 7.445000 0.580000 7.735000 0.625000 ;
  END
END sky130_fd_sc_hd__xor3_1
MACRO sky130_fd_sc_hd__xor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.965000 1.075000 8.375000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.145000 0.995000 7.315000 1.445000 ;
        RECT 7.145000 1.445000 7.725000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.320000 0.995000 2.955000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.660000 1.050000 0.925000 ;
        RECT 0.545000 0.925000 0.860000 1.440000 ;
        RECT 0.545000 1.440000 1.070000 2.045000 ;
        RECT 0.800000 0.350000 1.050000 0.660000 ;
        RECT 0.820000 2.045000 1.070000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.300000  0.085000 0.630000 0.465000 ;
      RECT 0.300000  2.215000 0.650000 2.635000 ;
      RECT 1.210000  0.995000 1.410000 1.325000 ;
      RECT 1.220000  0.085000 1.470000 0.525000 ;
      RECT 1.240000  0.695000 1.810000 0.865000 ;
      RECT 1.240000  0.865000 1.410000 0.995000 ;
      RECT 1.240000  1.325000 1.410000 1.875000 ;
      RECT 1.240000  1.875000 1.930000 2.045000 ;
      RECT 1.240000  2.215000 1.575000 2.635000 ;
      RECT 1.640000  0.255000 3.200000 0.425000 ;
      RECT 1.640000  0.425000 1.810000 0.695000 ;
      RECT 1.645000  1.535000 3.295000 1.705000 ;
      RECT 1.760000  2.045000 1.930000 2.235000 ;
      RECT 1.760000  2.235000 3.355000 2.405000 ;
      RECT 1.980000  0.595000 2.150000 1.535000 ;
      RECT 2.330000  1.895000 3.635000 2.065000 ;
      RECT 2.430000  0.655000 3.540000 0.825000 ;
      RECT 2.850000  0.425000 3.200000 0.455000 ;
      RECT 3.125000  0.995000 3.400000 1.325000 ;
      RECT 3.125000  1.325000 3.295000 1.535000 ;
      RECT 3.370000  0.255000 4.220000 0.425000 ;
      RECT 3.370000  0.425000 3.540000 0.655000 ;
      RECT 3.465000  1.525000 3.995000 1.695000 ;
      RECT 3.465000  1.695000 3.635000 1.895000 ;
      RECT 3.570000  2.235000 3.975000 2.405000 ;
      RECT 3.710000  0.595000 3.880000 1.375000 ;
      RECT 3.710000  1.375000 3.995000 1.525000 ;
      RECT 3.805000  1.895000 4.980000 2.065000 ;
      RECT 3.805000  2.065000 3.975000 2.235000 ;
      RECT 4.050000  0.425000 4.220000 1.035000 ;
      RECT 4.050000  1.035000 4.335000 1.205000 ;
      RECT 4.145000  2.235000 4.475000 2.635000 ;
      RECT 4.165000  1.205000 4.335000 1.895000 ;
      RECT 4.390000  0.085000 4.560000 0.865000 ;
      RECT 4.565000  1.445000 4.980000 1.715000 ;
      RECT 4.740000  0.415000 4.980000 1.445000 ;
      RECT 4.810000  2.065000 4.980000 2.275000 ;
      RECT 4.810000  2.275000 7.905000 2.445000 ;
      RECT 5.155000  0.265000 5.570000 0.485000 ;
      RECT 5.155000  0.485000 5.375000 0.595000 ;
      RECT 5.155000  0.595000 5.325000 2.105000 ;
      RECT 5.495000  0.720000 5.910000 0.825000 ;
      RECT 5.495000  0.825000 5.715000 0.890000 ;
      RECT 5.495000  0.890000 5.665000 2.275000 ;
      RECT 5.545000  0.655000 5.910000 0.720000 ;
      RECT 5.740000  0.320000 5.910000 0.655000 ;
      RECT 5.855000  1.445000 6.635000 1.615000 ;
      RECT 5.855000  1.615000 6.270000 2.045000 ;
      RECT 5.870000  0.995000 6.295000 1.270000 ;
      RECT 6.080000  0.630000 6.295000 0.995000 ;
      RECT 6.465000  0.255000 7.610000 0.425000 ;
      RECT 6.465000  0.425000 6.635000 1.445000 ;
      RECT 6.805000  0.595000 6.975000 1.935000 ;
      RECT 6.805000  1.935000 9.115000 2.105000 ;
      RECT 7.145000  0.425000 7.610000 0.465000 ;
      RECT 7.485000  0.730000 7.690000 0.945000 ;
      RECT 7.485000  0.945000 7.795000 1.275000 ;
      RECT 7.895000  1.495000 8.715000 1.705000 ;
      RECT 7.935000  0.295000 8.225000 0.735000 ;
      RECT 7.935000  0.735000 8.715000 0.750000 ;
      RECT 7.975000  0.750000 8.715000 0.905000 ;
      RECT 8.315000  2.275000 8.650000 2.635000 ;
      RECT 8.395000  0.085000 8.565000 0.565000 ;
      RECT 8.545000  0.905000 8.715000 0.995000 ;
      RECT 8.545000  0.995000 8.775000 1.325000 ;
      RECT 8.545000  1.325000 8.715000 1.495000 ;
      RECT 8.630000  1.875000 9.115000 1.935000 ;
      RECT 8.815000  0.255000 9.115000 0.585000 ;
      RECT 8.820000  2.105000 9.115000 2.465000 ;
      RECT 8.945000  0.585000 9.115000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  1.445000 3.995000 1.615000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  0.765000 4.915000 0.935000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  0.425000 5.375000 0.595000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  0.765000 6.295000 0.935000 ;
      RECT 6.125000  1.445000 6.295000 1.615000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  0.765000 7.675000 0.935000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  0.425000 8.135000 0.595000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
    LAYER met1 ;
      RECT 3.765000 1.415000 4.055000 1.460000 ;
      RECT 3.765000 1.460000 6.355000 1.600000 ;
      RECT 3.765000 1.600000 4.055000 1.645000 ;
      RECT 4.685000 0.735000 4.975000 0.780000 ;
      RECT 4.685000 0.780000 7.735000 0.920000 ;
      RECT 4.685000 0.920000 4.975000 0.965000 ;
      RECT 5.145000 0.395000 5.435000 0.440000 ;
      RECT 5.145000 0.440000 8.195000 0.580000 ;
      RECT 5.145000 0.580000 5.435000 0.625000 ;
      RECT 6.065000 0.735000 6.355000 0.780000 ;
      RECT 6.065000 0.920000 6.355000 0.965000 ;
      RECT 6.065000 1.415000 6.355000 1.460000 ;
      RECT 6.065000 1.600000 6.355000 1.645000 ;
      RECT 7.445000 0.735000 7.735000 0.780000 ;
      RECT 7.445000 0.920000 7.735000 0.965000 ;
      RECT 7.905000 0.395000 8.195000 0.440000 ;
      RECT 7.905000 0.580000 8.195000 0.625000 ;
  END
END sky130_fd_sc_hd__xor3_2
MACRO sky130_fd_sc_hd__xor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.525000 1.075000 8.935000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.705000 0.995000 7.875000 1.445000 ;
        RECT 7.705000 1.445000 8.285000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.880000 0.995000 3.515000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.350000 0.765000 0.660000 ;
        RECT 0.595000 0.660000 1.605000 0.830000 ;
        RECT 0.595000 0.830000 1.535000 0.925000 ;
        RECT 0.695000 1.440000 1.420000 1.455000 ;
        RECT 0.695000 1.455000 1.705000 2.045000 ;
        RECT 0.695000 2.045000 0.865000 2.465000 ;
        RECT 1.105000 0.925000 1.420000 1.440000 ;
        RECT 1.435000 0.350000 1.605000 0.660000 ;
        RECT 1.535000 2.045000 1.705000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.120000 0.085000 ;
        RECT 0.175000  0.085000  0.345000 0.545000 ;
        RECT 0.935000  0.085000  1.265000 0.465000 ;
        RECT 1.855000  0.085000  2.025000 0.525000 ;
        RECT 4.950000  0.085000  5.120000 0.885000 ;
        RECT 8.995000  0.085000  9.165000 0.565000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
        RECT 7.965000 -0.085000 8.135000 0.085000 ;
        RECT 8.425000 -0.085000 8.595000 0.085000 ;
        RECT 8.885000 -0.085000 9.055000 0.085000 ;
        RECT 9.345000 -0.085000 9.515000 0.085000 ;
        RECT 9.805000 -0.085000 9.975000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.235000 -0.085000 0.405000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 10.120000 2.805000 ;
        RECT 0.275000 2.135000  0.445000 2.635000 ;
        RECT 1.035000 2.215000  1.365000 2.635000 ;
        RECT 1.875000 2.215000  2.205000 2.635000 ;
        RECT 4.705000 2.235000  5.035000 2.635000 ;
        RECT 8.915000 2.275000  9.245000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
        RECT 8.425000 2.635000 8.595000 2.805000 ;
        RECT 8.885000 2.635000 9.055000 2.805000 ;
        RECT 9.345000 2.635000 9.515000 2.805000 ;
        RECT 9.805000 2.635000 9.975000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.820000 0.965000 2.045000 1.325000 ;
      RECT 1.875000 0.695000 2.365000 0.865000 ;
      RECT 1.875000 0.865000 2.045000 0.965000 ;
      RECT 1.875000 1.325000 2.045000 1.875000 ;
      RECT 1.875000 1.875000 2.545000 2.045000 ;
      RECT 2.195000 0.255000 3.760000 0.425000 ;
      RECT 2.195000 0.425000 2.365000 0.695000 ;
      RECT 2.370000 1.535000 3.855000 1.705000 ;
      RECT 2.375000 2.045000 2.545000 2.235000 ;
      RECT 2.375000 2.235000 3.915000 2.405000 ;
      RECT 2.540000 0.595000 2.710000 1.535000 ;
      RECT 2.890000 1.895000 4.195000 2.065000 ;
      RECT 2.990000 0.655000 4.100000 0.825000 ;
      RECT 3.410000 0.425000 3.760000 0.455000 ;
      RECT 3.685000 0.995000 4.055000 1.325000 ;
      RECT 3.685000 1.325000 3.855000 1.535000 ;
      RECT 3.930000 0.255000 4.780000 0.425000 ;
      RECT 3.930000 0.425000 4.100000 0.655000 ;
      RECT 4.025000 1.525000 4.555000 1.695000 ;
      RECT 4.025000 1.695000 4.195000 1.895000 ;
      RECT 4.130000 2.235000 4.535000 2.405000 ;
      RECT 4.270000 0.595000 4.440000 1.375000 ;
      RECT 4.270000 1.375000 4.555000 1.525000 ;
      RECT 4.365000 1.895000 5.540000 2.065000 ;
      RECT 4.365000 2.065000 4.535000 2.235000 ;
      RECT 4.610000 0.425000 4.780000 1.035000 ;
      RECT 4.610000 1.035000 4.865000 1.040000 ;
      RECT 4.610000 1.040000 4.880000 1.045000 ;
      RECT 4.610000 1.045000 4.890000 1.050000 ;
      RECT 4.610000 1.050000 4.895000 1.205000 ;
      RECT 4.725000 1.205000 4.895000 1.895000 ;
      RECT 5.125000 1.445000 5.540000 1.715000 ;
      RECT 5.300000 0.415000 5.540000 1.445000 ;
      RECT 5.370000 2.065000 5.540000 2.275000 ;
      RECT 5.370000 2.275000 8.465000 2.445000 ;
      RECT 5.715000 0.265000 6.130000 0.485000 ;
      RECT 5.715000 0.485000 5.935000 0.595000 ;
      RECT 5.715000 0.595000 5.885000 2.105000 ;
      RECT 6.075000 0.720000 6.470000 0.825000 ;
      RECT 6.075000 0.825000 6.275000 0.890000 ;
      RECT 6.075000 0.890000 6.245000 2.275000 ;
      RECT 6.105000 0.655000 6.470000 0.720000 ;
      RECT 6.300000 0.320000 6.470000 0.655000 ;
      RECT 6.415000 1.445000 7.195000 1.615000 ;
      RECT 6.415000 1.615000 6.830000 2.045000 ;
      RECT 6.430000 0.995000 6.855000 1.270000 ;
      RECT 6.640000 0.630000 6.855000 0.995000 ;
      RECT 7.025000 0.255000 8.170000 0.425000 ;
      RECT 7.025000 0.425000 7.195000 1.445000 ;
      RECT 7.365000 0.595000 7.535000 1.935000 ;
      RECT 7.365000 1.935000 9.675000 2.105000 ;
      RECT 7.705000 0.425000 8.170000 0.465000 ;
      RECT 8.045000 0.730000 8.250000 0.945000 ;
      RECT 8.045000 0.945000 8.355000 1.275000 ;
      RECT 8.455000 1.495000 9.275000 1.705000 ;
      RECT 8.495000 0.295000 8.785000 0.735000 ;
      RECT 8.495000 0.735000 9.275000 0.750000 ;
      RECT 8.535000 0.750000 9.275000 0.905000 ;
      RECT 9.105000 0.905000 9.275000 0.995000 ;
      RECT 9.105000 0.995000 9.335000 1.325000 ;
      RECT 9.105000 1.325000 9.275000 1.495000 ;
      RECT 9.190000 1.875000 9.675000 1.935000 ;
      RECT 9.415000 0.255000 9.675000 0.585000 ;
      RECT 9.415000 2.105000 9.675000 2.465000 ;
      RECT 9.505000 0.585000 9.675000 1.875000 ;
    LAYER mcon ;
      RECT 4.385000 1.445000 4.555000 1.615000 ;
      RECT 5.305000 0.765000 5.475000 0.935000 ;
      RECT 5.765000 0.425000 5.935000 0.595000 ;
      RECT 6.685000 0.765000 6.855000 0.935000 ;
      RECT 6.685000 1.445000 6.855000 1.615000 ;
      RECT 8.065000 0.765000 8.235000 0.935000 ;
      RECT 8.525000 0.425000 8.695000 0.595000 ;
    LAYER met1 ;
      RECT 4.325000 1.415000 4.615000 1.460000 ;
      RECT 4.325000 1.460000 6.915000 1.600000 ;
      RECT 4.325000 1.600000 4.615000 1.645000 ;
      RECT 5.245000 0.735000 5.535000 0.780000 ;
      RECT 5.245000 0.780000 8.295000 0.920000 ;
      RECT 5.245000 0.920000 5.535000 0.965000 ;
      RECT 5.705000 0.395000 5.995000 0.440000 ;
      RECT 5.705000 0.440000 8.755000 0.580000 ;
      RECT 5.705000 0.580000 5.995000 0.625000 ;
      RECT 6.625000 0.735000 6.915000 0.780000 ;
      RECT 6.625000 0.920000 6.915000 0.965000 ;
      RECT 6.625000 1.415000 6.915000 1.460000 ;
      RECT 6.625000 1.600000 6.915000 1.645000 ;
      RECT 8.005000 0.735000 8.295000 0.780000 ;
      RECT 8.005000 0.920000 8.295000 0.965000 ;
      RECT 8.465000 0.395000 8.755000 0.440000 ;
      RECT 8.465000 0.580000 8.755000 0.625000 ;
  END
END sky130_fd_sc_hd__xor3_4
MACRO qspim_top
  CLASS BLOCK ;
  FOREIGN qspim_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 650.000 ;
  PIN mclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 0.720 4.000 1.320 ;
    END
  END mclk
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2.080 4.000 2.680 ;
    END
  END rst_n
  PIN spi_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 211.520 404.000 212.120 ;
    END
  END spi_clk
  PIN spi_csn0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 212.880 404.000 213.480 ;
    END
  END spi_csn0
  PIN spi_debug[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 0.720 404.000 1.320 ;
    END
  END spi_debug[0]
  PIN spi_debug[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 14.320 404.000 14.920 ;
    END
  END spi_debug[10]
  PIN spi_debug[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 15.680 404.000 16.280 ;
    END
  END spi_debug[11]
  PIN spi_debug[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 17.040 404.000 17.640 ;
    END
  END spi_debug[12]
  PIN spi_debug[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 18.400 404.000 19.000 ;
    END
  END spi_debug[13]
  PIN spi_debug[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 19.760 404.000 20.360 ;
    END
  END spi_debug[14]
  PIN spi_debug[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 21.120 404.000 21.720 ;
    END
  END spi_debug[15]
  PIN spi_debug[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 22.480 404.000 23.080 ;
    END
  END spi_debug[16]
  PIN spi_debug[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 23.840 404.000 24.440 ;
    END
  END spi_debug[17]
  PIN spi_debug[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 25.200 404.000 25.800 ;
    END
  END spi_debug[18]
  PIN spi_debug[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 26.560 404.000 27.160 ;
    END
  END spi_debug[19]
  PIN spi_debug[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 2.080 404.000 2.680 ;
    END
  END spi_debug[1]
  PIN spi_debug[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 27.920 404.000 28.520 ;
    END
  END spi_debug[20]
  PIN spi_debug[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 29.280 404.000 29.880 ;
    END
  END spi_debug[21]
  PIN spi_debug[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 30.640 404.000 31.240 ;
    END
  END spi_debug[22]
  PIN spi_debug[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 32.000 404.000 32.600 ;
    END
  END spi_debug[23]
  PIN spi_debug[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 33.360 404.000 33.960 ;
    END
  END spi_debug[24]
  PIN spi_debug[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 34.720 404.000 35.320 ;
    END
  END spi_debug[25]
  PIN spi_debug[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 36.080 404.000 36.680 ;
    END
  END spi_debug[26]
  PIN spi_debug[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 37.440 404.000 38.040 ;
    END
  END spi_debug[27]
  PIN spi_debug[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 38.800 404.000 39.400 ;
    END
  END spi_debug[28]
  PIN spi_debug[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 40.160 404.000 40.760 ;
    END
  END spi_debug[29]
  PIN spi_debug[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 3.440 404.000 4.040 ;
    END
  END spi_debug[2]
  PIN spi_debug[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 41.520 404.000 42.120 ;
    END
  END spi_debug[30]
  PIN spi_debug[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 42.880 404.000 43.480 ;
    END
  END spi_debug[31]
  PIN spi_debug[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 4.800 404.000 5.400 ;
    END
  END spi_debug[3]
  PIN spi_debug[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 6.160 404.000 6.760 ;
    END
  END spi_debug[4]
  PIN spi_debug[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 7.520 404.000 8.120 ;
    END
  END spi_debug[5]
  PIN spi_debug[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 8.880 404.000 9.480 ;
    END
  END spi_debug[6]
  PIN spi_debug[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 10.240 404.000 10.840 ;
    END
  END spi_debug[7]
  PIN spi_debug[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 11.600 404.000 12.200 ;
    END
  END spi_debug[8]
  PIN spi_debug[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 12.960 404.000 13.560 ;
    END
  END spi_debug[9]
  PIN spi_oen[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 218.320 404.000 218.920 ;
    END
  END spi_oen[0]
  PIN spi_oen[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 216.960 404.000 217.560 ;
    END
  END spi_oen[1]
  PIN spi_oen[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 215.600 404.000 216.200 ;
    END
  END spi_oen[2]
  PIN spi_oen[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 214.240 404.000 214.840 ;
    END
  END spi_oen[3]
  PIN spi_sdi[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 204.720 404.000 205.320 ;
    END
  END spi_sdi[0]
  PIN spi_sdi[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 203.360 404.000 203.960 ;
    END
  END spi_sdi[1]
  PIN spi_sdi[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 202.000 404.000 202.600 ;
    END
  END spi_sdi[2]
  PIN spi_sdi[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 200.640 404.000 201.240 ;
    END
  END spi_sdi[3]
  PIN spi_sdo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 210.160 404.000 210.760 ;
    END
  END spi_sdo[0]
  PIN spi_sdo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 208.800 404.000 209.400 ;
    END
  END spi_sdo[1]
  PIN spi_sdo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 207.440 404.000 208.040 ;
    END
  END spi_sdo[2]
  PIN spi_sdo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 206.080 404.000 206.680 ;
    END
  END spi_sdo[3]
  PIN wbd_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 -4.000 94.670 4.000 ;
    END
  END wbd_ack_o
  PIN wbd_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 -4.000 31.190 4.000 ;
    END
  END wbd_adr_i[0]
  PIN wbd_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 -4.000 21.990 4.000 ;
    END
  END wbd_adr_i[10]
  PIN wbd_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 -4.000 21.070 4.000 ;
    END
  END wbd_adr_i[11]
  PIN wbd_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 -4.000 20.150 4.000 ;
    END
  END wbd_adr_i[12]
  PIN wbd_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 -4.000 19.230 4.000 ;
    END
  END wbd_adr_i[13]
  PIN wbd_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 -4.000 18.310 4.000 ;
    END
  END wbd_adr_i[14]
  PIN wbd_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 -4.000 17.390 4.000 ;
    END
  END wbd_adr_i[15]
  PIN wbd_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 -4.000 16.470 4.000 ;
    END
  END wbd_adr_i[16]
  PIN wbd_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 -4.000 15.550 4.000 ;
    END
  END wbd_adr_i[17]
  PIN wbd_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 -4.000 14.630 4.000 ;
    END
  END wbd_adr_i[18]
  PIN wbd_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 -4.000 13.710 4.000 ;
    END
  END wbd_adr_i[19]
  PIN wbd_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 -4.000 30.270 4.000 ;
    END
  END wbd_adr_i[1]
  PIN wbd_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 -4.000 12.790 4.000 ;
    END
  END wbd_adr_i[20]
  PIN wbd_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 -4.000 11.870 4.000 ;
    END
  END wbd_adr_i[21]
  PIN wbd_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 -4.000 10.950 4.000 ;
    END
  END wbd_adr_i[22]
  PIN wbd_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 -4.000 10.030 4.000 ;
    END
  END wbd_adr_i[23]
  PIN wbd_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 -4.000 9.110 4.000 ;
    END
  END wbd_adr_i[24]
  PIN wbd_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 -4.000 8.190 4.000 ;
    END
  END wbd_adr_i[25]
  PIN wbd_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 -4.000 7.270 4.000 ;
    END
  END wbd_adr_i[26]
  PIN wbd_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 -4.000 6.350 4.000 ;
    END
  END wbd_adr_i[27]
  PIN wbd_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 -4.000 5.430 4.000 ;
    END
  END wbd_adr_i[28]
  PIN wbd_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 -4.000 4.510 4.000 ;
    END
  END wbd_adr_i[29]
  PIN wbd_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 -4.000 29.350 4.000 ;
    END
  END wbd_adr_i[2]
  PIN wbd_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 -4.000 3.590 4.000 ;
    END
  END wbd_adr_i[30]
  PIN wbd_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 -4.000 2.670 4.000 ;
    END
  END wbd_adr_i[31]
  PIN wbd_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 -4.000 28.430 4.000 ;
    END
  END wbd_adr_i[3]
  PIN wbd_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 -4.000 27.510 4.000 ;
    END
  END wbd_adr_i[4]
  PIN wbd_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 -4.000 26.590 4.000 ;
    END
  END wbd_adr_i[5]
  PIN wbd_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 -4.000 25.670 4.000 ;
    END
  END wbd_adr_i[6]
  PIN wbd_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 -4.000 24.750 4.000 ;
    END
  END wbd_adr_i[7]
  PIN wbd_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 -4.000 23.830 4.000 ;
    END
  END wbd_adr_i[8]
  PIN wbd_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 -4.000 22.910 4.000 ;
    END
  END wbd_adr_i[9]
  PIN wbd_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 -4.000 64.310 4.000 ;
    END
  END wbd_dat_i[0]
  PIN wbd_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 -4.000 55.110 4.000 ;
    END
  END wbd_dat_i[10]
  PIN wbd_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 -4.000 54.190 4.000 ;
    END
  END wbd_dat_i[11]
  PIN wbd_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 -4.000 53.270 4.000 ;
    END
  END wbd_dat_i[12]
  PIN wbd_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 -4.000 52.350 4.000 ;
    END
  END wbd_dat_i[13]
  PIN wbd_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 -4.000 51.430 4.000 ;
    END
  END wbd_dat_i[14]
  PIN wbd_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 -4.000 50.510 4.000 ;
    END
  END wbd_dat_i[15]
  PIN wbd_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 -4.000 49.590 4.000 ;
    END
  END wbd_dat_i[16]
  PIN wbd_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 -4.000 48.670 4.000 ;
    END
  END wbd_dat_i[17]
  PIN wbd_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 -4.000 47.750 4.000 ;
    END
  END wbd_dat_i[18]
  PIN wbd_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 -4.000 46.830 4.000 ;
    END
  END wbd_dat_i[19]
  PIN wbd_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 -4.000 63.390 4.000 ;
    END
  END wbd_dat_i[1]
  PIN wbd_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 -4.000 45.910 4.000 ;
    END
  END wbd_dat_i[20]
  PIN wbd_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 -4.000 44.990 4.000 ;
    END
  END wbd_dat_i[21]
  PIN wbd_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 -4.000 44.070 4.000 ;
    END
  END wbd_dat_i[22]
  PIN wbd_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 -4.000 43.150 4.000 ;
    END
  END wbd_dat_i[23]
  PIN wbd_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 -4.000 42.230 4.000 ;
    END
  END wbd_dat_i[24]
  PIN wbd_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 -4.000 41.310 4.000 ;
    END
  END wbd_dat_i[25]
  PIN wbd_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 -4.000 40.390 4.000 ;
    END
  END wbd_dat_i[26]
  PIN wbd_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 -4.000 39.470 4.000 ;
    END
  END wbd_dat_i[27]
  PIN wbd_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 -4.000 38.550 4.000 ;
    END
  END wbd_dat_i[28]
  PIN wbd_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 -4.000 37.630 4.000 ;
    END
  END wbd_dat_i[29]
  PIN wbd_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 -4.000 62.470 4.000 ;
    END
  END wbd_dat_i[2]
  PIN wbd_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 -4.000 36.710 4.000 ;
    END
  END wbd_dat_i[30]
  PIN wbd_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 -4.000 35.790 4.000 ;
    END
  END wbd_dat_i[31]
  PIN wbd_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 -4.000 61.550 4.000 ;
    END
  END wbd_dat_i[3]
  PIN wbd_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 -4.000 60.630 4.000 ;
    END
  END wbd_dat_i[4]
  PIN wbd_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 -4.000 59.710 4.000 ;
    END
  END wbd_dat_i[5]
  PIN wbd_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 -4.000 58.790 4.000 ;
    END
  END wbd_dat_i[6]
  PIN wbd_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 -4.000 57.870 4.000 ;
    END
  END wbd_dat_i[7]
  PIN wbd_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 -4.000 56.950 4.000 ;
    END
  END wbd_dat_i[8]
  PIN wbd_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 -4.000 56.030 4.000 ;
    END
  END wbd_dat_i[9]
  PIN wbd_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 -4.000 93.750 4.000 ;
    END
  END wbd_dat_o[0]
  PIN wbd_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 -4.000 84.550 4.000 ;
    END
  END wbd_dat_o[10]
  PIN wbd_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 -4.000 83.630 4.000 ;
    END
  END wbd_dat_o[11]
  PIN wbd_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 -4.000 82.710 4.000 ;
    END
  END wbd_dat_o[12]
  PIN wbd_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 -4.000 81.790 4.000 ;
    END
  END wbd_dat_o[13]
  PIN wbd_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 -4.000 80.870 4.000 ;
    END
  END wbd_dat_o[14]
  PIN wbd_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 -4.000 79.950 4.000 ;
    END
  END wbd_dat_o[15]
  PIN wbd_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 -4.000 79.030 4.000 ;
    END
  END wbd_dat_o[16]
  PIN wbd_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 -4.000 78.110 4.000 ;
    END
  END wbd_dat_o[17]
  PIN wbd_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 -4.000 77.190 4.000 ;
    END
  END wbd_dat_o[18]
  PIN wbd_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 -4.000 76.270 4.000 ;
    END
  END wbd_dat_o[19]
  PIN wbd_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 -4.000 92.830 4.000 ;
    END
  END wbd_dat_o[1]
  PIN wbd_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 -4.000 75.350 4.000 ;
    END
  END wbd_dat_o[20]
  PIN wbd_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 -4.000 74.430 4.000 ;
    END
  END wbd_dat_o[21]
  PIN wbd_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 -4.000 73.510 4.000 ;
    END
  END wbd_dat_o[22]
  PIN wbd_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 -4.000 72.590 4.000 ;
    END
  END wbd_dat_o[23]
  PIN wbd_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 -4.000 71.670 4.000 ;
    END
  END wbd_dat_o[24]
  PIN wbd_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 -4.000 70.750 4.000 ;
    END
  END wbd_dat_o[25]
  PIN wbd_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 -4.000 69.830 4.000 ;
    END
  END wbd_dat_o[26]
  PIN wbd_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 -4.000 68.910 4.000 ;
    END
  END wbd_dat_o[27]
  PIN wbd_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 -4.000 67.990 4.000 ;
    END
  END wbd_dat_o[28]
  PIN wbd_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 -4.000 67.070 4.000 ;
    END
  END wbd_dat_o[29]
  PIN wbd_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 -4.000 91.910 4.000 ;
    END
  END wbd_dat_o[2]
  PIN wbd_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 -4.000 66.150 4.000 ;
    END
  END wbd_dat_o[30]
  PIN wbd_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 -4.000 65.230 4.000 ;
    END
  END wbd_dat_o[31]
  PIN wbd_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 -4.000 90.990 4.000 ;
    END
  END wbd_dat_o[3]
  PIN wbd_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 -4.000 90.070 4.000 ;
    END
  END wbd_dat_o[4]
  PIN wbd_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 -4.000 89.150 4.000 ;
    END
  END wbd_dat_o[5]
  PIN wbd_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 -4.000 88.230 4.000 ;
    END
  END wbd_dat_o[6]
  PIN wbd_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 -4.000 87.310 4.000 ;
    END
  END wbd_dat_o[7]
  PIN wbd_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 -4.000 86.390 4.000 ;
    END
  END wbd_dat_o[8]
  PIN wbd_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 -4.000 85.470 4.000 ;
    END
  END wbd_dat_o[9]
  PIN wbd_err_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 -4.000 95.590 4.000 ;
    END
  END wbd_err_o
  PIN wbd_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 -4.000 34.870 4.000 ;
    END
  END wbd_sel_i[0]
  PIN wbd_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 -4.000 33.950 4.000 ;
    END
  END wbd_sel_i[1]
  PIN wbd_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 -4.000 33.030 4.000 ;
    END
  END wbd_sel_i[2]
  PIN wbd_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 -4.000 32.110 4.000 ;
    END
  END wbd_sel_i[3]
  PIN wbd_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 -4.000 0.830 4.000 ;
    END
  END wbd_stb_i
  PIN wbd_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 -4.000 1.750 4.000 ;
    END
  END wbd_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 319.340 10.640 324.340 636.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 219.340 10.640 224.340 636.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 119.340 10.640 124.340 636.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.340 10.640 24.340 636.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 369.340 10.640 374.340 636.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 269.340 10.640 274.340 636.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 169.340 10.640 174.340 636.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 69.340 10.640 74.340 636.720 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 394.995 636.565 ;
      LAYER met1 ;
        RECT 0.530 3.100 395.055 636.720 ;
      LAYER met2 ;
        RECT 0.560 4.280 392.290 636.720 ;
        RECT 1.110 0.835 1.190 4.280 ;
        RECT 2.030 0.835 2.110 4.280 ;
        RECT 2.950 0.835 3.030 4.280 ;
        RECT 3.870 0.835 3.950 4.280 ;
        RECT 4.790 0.835 4.870 4.280 ;
        RECT 5.710 0.835 5.790 4.280 ;
        RECT 6.630 0.835 6.710 4.280 ;
        RECT 7.550 0.835 7.630 4.280 ;
        RECT 8.470 0.835 8.550 4.280 ;
        RECT 9.390 0.835 9.470 4.280 ;
        RECT 10.310 0.835 10.390 4.280 ;
        RECT 11.230 0.835 11.310 4.280 ;
        RECT 12.150 0.835 12.230 4.280 ;
        RECT 13.070 0.835 13.150 4.280 ;
        RECT 13.990 0.835 14.070 4.280 ;
        RECT 14.910 0.835 14.990 4.280 ;
        RECT 15.830 0.835 15.910 4.280 ;
        RECT 16.750 0.835 16.830 4.280 ;
        RECT 17.670 0.835 17.750 4.280 ;
        RECT 18.590 0.835 18.670 4.280 ;
        RECT 19.510 0.835 19.590 4.280 ;
        RECT 20.430 0.835 20.510 4.280 ;
        RECT 21.350 0.835 21.430 4.280 ;
        RECT 22.270 0.835 22.350 4.280 ;
        RECT 23.190 0.835 23.270 4.280 ;
        RECT 24.110 0.835 24.190 4.280 ;
        RECT 25.030 0.835 25.110 4.280 ;
        RECT 25.950 0.835 26.030 4.280 ;
        RECT 26.870 0.835 26.950 4.280 ;
        RECT 27.790 0.835 27.870 4.280 ;
        RECT 28.710 0.835 28.790 4.280 ;
        RECT 29.630 0.835 29.710 4.280 ;
        RECT 30.550 0.835 30.630 4.280 ;
        RECT 31.470 0.835 31.550 4.280 ;
        RECT 32.390 0.835 32.470 4.280 ;
        RECT 33.310 0.835 33.390 4.280 ;
        RECT 34.230 0.835 34.310 4.280 ;
        RECT 35.150 0.835 35.230 4.280 ;
        RECT 36.070 0.835 36.150 4.280 ;
        RECT 36.990 0.835 37.070 4.280 ;
        RECT 37.910 0.835 37.990 4.280 ;
        RECT 38.830 0.835 38.910 4.280 ;
        RECT 39.750 0.835 39.830 4.280 ;
        RECT 40.670 0.835 40.750 4.280 ;
        RECT 41.590 0.835 41.670 4.280 ;
        RECT 42.510 0.835 42.590 4.280 ;
        RECT 43.430 0.835 43.510 4.280 ;
        RECT 44.350 0.835 44.430 4.280 ;
        RECT 45.270 0.835 45.350 4.280 ;
        RECT 46.190 0.835 46.270 4.280 ;
        RECT 47.110 0.835 47.190 4.280 ;
        RECT 48.030 0.835 48.110 4.280 ;
        RECT 48.950 0.835 49.030 4.280 ;
        RECT 49.870 0.835 49.950 4.280 ;
        RECT 50.790 0.835 50.870 4.280 ;
        RECT 51.710 0.835 51.790 4.280 ;
        RECT 52.630 0.835 52.710 4.280 ;
        RECT 53.550 0.835 53.630 4.280 ;
        RECT 54.470 0.835 54.550 4.280 ;
        RECT 55.390 0.835 55.470 4.280 ;
        RECT 56.310 0.835 56.390 4.280 ;
        RECT 57.230 0.835 57.310 4.280 ;
        RECT 58.150 0.835 58.230 4.280 ;
        RECT 59.070 0.835 59.150 4.280 ;
        RECT 59.990 0.835 60.070 4.280 ;
        RECT 60.910 0.835 60.990 4.280 ;
        RECT 61.830 0.835 61.910 4.280 ;
        RECT 62.750 0.835 62.830 4.280 ;
        RECT 63.670 0.835 63.750 4.280 ;
        RECT 64.590 0.835 64.670 4.280 ;
        RECT 65.510 0.835 65.590 4.280 ;
        RECT 66.430 0.835 66.510 4.280 ;
        RECT 67.350 0.835 67.430 4.280 ;
        RECT 68.270 0.835 68.350 4.280 ;
        RECT 69.190 0.835 69.270 4.280 ;
        RECT 70.110 0.835 70.190 4.280 ;
        RECT 71.030 0.835 71.110 4.280 ;
        RECT 71.950 0.835 72.030 4.280 ;
        RECT 72.870 0.835 72.950 4.280 ;
        RECT 73.790 0.835 73.870 4.280 ;
        RECT 74.710 0.835 74.790 4.280 ;
        RECT 75.630 0.835 75.710 4.280 ;
        RECT 76.550 0.835 76.630 4.280 ;
        RECT 77.470 0.835 77.550 4.280 ;
        RECT 78.390 0.835 78.470 4.280 ;
        RECT 79.310 0.835 79.390 4.280 ;
        RECT 80.230 0.835 80.310 4.280 ;
        RECT 81.150 0.835 81.230 4.280 ;
        RECT 82.070 0.835 82.150 4.280 ;
        RECT 82.990 0.835 83.070 4.280 ;
        RECT 83.910 0.835 83.990 4.280 ;
        RECT 84.830 0.835 84.910 4.280 ;
        RECT 85.750 0.835 85.830 4.280 ;
        RECT 86.670 0.835 86.750 4.280 ;
        RECT 87.590 0.835 87.670 4.280 ;
        RECT 88.510 0.835 88.590 4.280 ;
        RECT 89.430 0.835 89.510 4.280 ;
        RECT 90.350 0.835 90.430 4.280 ;
        RECT 91.270 0.835 91.350 4.280 ;
        RECT 92.190 0.835 92.270 4.280 ;
        RECT 93.110 0.835 93.190 4.280 ;
        RECT 94.030 0.835 94.110 4.280 ;
        RECT 94.950 0.835 95.030 4.280 ;
        RECT 95.870 0.835 392.290 4.280 ;
      LAYER met3 ;
        RECT 4.000 219.320 396.000 636.645 ;
        RECT 4.000 200.240 395.600 219.320 ;
        RECT 4.000 43.880 396.000 200.240 ;
        RECT 4.000 3.080 395.600 43.880 ;
        RECT 4.400 0.855 395.600 3.080 ;
  END
END qspim_top
MACRO pinmux
  CLASS BLOCK ;
  FOREIGN pinmux ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN digital_io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 0.720 504.000 1.320 ;
    END
  END digital_io_in[0]
  PIN digital_io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 82.320 504.000 82.920 ;
    END
  END digital_io_in[10]
  PIN digital_io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 90.480 504.000 91.080 ;
    END
  END digital_io_in[11]
  PIN digital_io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 98.640 504.000 99.240 ;
    END
  END digital_io_in[12]
  PIN digital_io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 106.800 504.000 107.400 ;
    END
  END digital_io_in[13]
  PIN digital_io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 114.960 504.000 115.560 ;
    END
  END digital_io_in[14]
  PIN digital_io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 496.000 322.830 504.000 ;
    END
  END digital_io_in[15]
  PIN digital_io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 496.000 320.070 504.000 ;
    END
  END digital_io_in[16]
  PIN digital_io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 496.000 317.310 504.000 ;
    END
  END digital_io_in[17]
  PIN digital_io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 496.000 314.550 504.000 ;
    END
  END digital_io_in[18]
  PIN digital_io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 496.000 311.790 504.000 ;
    END
  END digital_io_in[19]
  PIN digital_io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 8.880 504.000 9.480 ;
    END
  END digital_io_in[1]
  PIN digital_io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 496.000 309.030 504.000 ;
    END
  END digital_io_in[20]
  PIN digital_io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 496.000 306.270 504.000 ;
    END
  END digital_io_in[21]
  PIN digital_io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 496.000 303.510 504.000 ;
    END
  END digital_io_in[22]
  PIN digital_io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 496.000 300.750 504.000 ;
    END
  END digital_io_in[23]
  PIN digital_io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 218.320 4.000 218.920 ;
    END
  END digital_io_in[24]
  PIN digital_io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 214.240 4.000 214.840 ;
    END
  END digital_io_in[25]
  PIN digital_io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 210.160 4.000 210.760 ;
    END
  END digital_io_in[26]
  PIN digital_io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 206.080 4.000 206.680 ;
    END
  END digital_io_in[27]
  PIN digital_io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 202.000 4.000 202.600 ;
    END
  END digital_io_in[28]
  PIN digital_io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 55.120 4.000 55.720 ;
    END
  END digital_io_in[29]
  PIN digital_io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 17.040 504.000 17.640 ;
    END
  END digital_io_in[2]
  PIN digital_io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 51.040 4.000 51.640 ;
    END
  END digital_io_in[30]
  PIN digital_io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 46.960 4.000 47.560 ;
    END
  END digital_io_in[31]
  PIN digital_io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 42.880 4.000 43.480 ;
    END
  END digital_io_in[32]
  PIN digital_io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 38.800 4.000 39.400 ;
    END
  END digital_io_in[33]
  PIN digital_io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 34.720 4.000 35.320 ;
    END
  END digital_io_in[34]
  PIN digital_io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 30.640 4.000 31.240 ;
    END
  END digital_io_in[35]
  PIN digital_io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 26.560 4.000 27.160 ;
    END
  END digital_io_in[36]
  PIN digital_io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 22.480 4.000 23.080 ;
    END
  END digital_io_in[37]
  PIN digital_io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 25.200 504.000 25.800 ;
    END
  END digital_io_in[3]
  PIN digital_io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 33.360 504.000 33.960 ;
    END
  END digital_io_in[4]
  PIN digital_io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 41.520 504.000 42.120 ;
    END
  END digital_io_in[5]
  PIN digital_io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 49.680 504.000 50.280 ;
    END
  END digital_io_in[6]
  PIN digital_io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 57.840 504.000 58.440 ;
    END
  END digital_io_in[7]
  PIN digital_io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 66.000 504.000 66.600 ;
    END
  END digital_io_in[8]
  PIN digital_io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 74.160 504.000 74.760 ;
    END
  END digital_io_in[9]
  PIN digital_io_oen[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 6.160 504.000 6.760 ;
    END
  END digital_io_oen[0]
  PIN digital_io_oen[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 87.760 504.000 88.360 ;
    END
  END digital_io_oen[10]
  PIN digital_io_oen[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 95.920 504.000 96.520 ;
    END
  END digital_io_oen[11]
  PIN digital_io_oen[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 104.080 504.000 104.680 ;
    END
  END digital_io_oen[12]
  PIN digital_io_oen[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 112.240 504.000 112.840 ;
    END
  END digital_io_oen[13]
  PIN digital_io_oen[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 120.400 504.000 121.000 ;
    END
  END digital_io_oen[14]
  PIN digital_io_oen[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 496.000 324.670 504.000 ;
    END
  END digital_io_oen[15]
  PIN digital_io_oen[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 496.000 321.910 504.000 ;
    END
  END digital_io_oen[16]
  PIN digital_io_oen[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 496.000 319.150 504.000 ;
    END
  END digital_io_oen[17]
  PIN digital_io_oen[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 496.000 316.390 504.000 ;
    END
  END digital_io_oen[18]
  PIN digital_io_oen[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 496.000 313.630 504.000 ;
    END
  END digital_io_oen[19]
  PIN digital_io_oen[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 14.320 504.000 14.920 ;
    END
  END digital_io_oen[1]
  PIN digital_io_oen[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 496.000 310.870 504.000 ;
    END
  END digital_io_oen[20]
  PIN digital_io_oen[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 496.000 308.110 504.000 ;
    END
  END digital_io_oen[21]
  PIN digital_io_oen[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 496.000 305.350 504.000 ;
    END
  END digital_io_oen[22]
  PIN digital_io_oen[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 496.000 302.590 504.000 ;
    END
  END digital_io_oen[23]
  PIN digital_io_oen[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 215.600 4.000 216.200 ;
    END
  END digital_io_oen[24]
  PIN digital_io_oen[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 211.520 4.000 212.120 ;
    END
  END digital_io_oen[25]
  PIN digital_io_oen[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 207.440 4.000 208.040 ;
    END
  END digital_io_oen[26]
  PIN digital_io_oen[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 203.360 4.000 203.960 ;
    END
  END digital_io_oen[27]
  PIN digital_io_oen[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 56.480 4.000 57.080 ;
    END
  END digital_io_oen[28]
  PIN digital_io_oen[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 52.400 4.000 53.000 ;
    END
  END digital_io_oen[29]
  PIN digital_io_oen[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 22.480 504.000 23.080 ;
    END
  END digital_io_oen[2]
  PIN digital_io_oen[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 48.320 4.000 48.920 ;
    END
  END digital_io_oen[30]
  PIN digital_io_oen[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 44.240 4.000 44.840 ;
    END
  END digital_io_oen[31]
  PIN digital_io_oen[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 40.160 4.000 40.760 ;
    END
  END digital_io_oen[32]
  PIN digital_io_oen[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 36.080 4.000 36.680 ;
    END
  END digital_io_oen[33]
  PIN digital_io_oen[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 32.000 4.000 32.600 ;
    END
  END digital_io_oen[34]
  PIN digital_io_oen[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 27.920 4.000 28.520 ;
    END
  END digital_io_oen[35]
  PIN digital_io_oen[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 23.840 4.000 24.440 ;
    END
  END digital_io_oen[36]
  PIN digital_io_oen[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 19.760 4.000 20.360 ;
    END
  END digital_io_oen[37]
  PIN digital_io_oen[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 30.640 504.000 31.240 ;
    END
  END digital_io_oen[3]
  PIN digital_io_oen[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 38.800 504.000 39.400 ;
    END
  END digital_io_oen[4]
  PIN digital_io_oen[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 46.960 504.000 47.560 ;
    END
  END digital_io_oen[5]
  PIN digital_io_oen[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 55.120 504.000 55.720 ;
    END
  END digital_io_oen[6]
  PIN digital_io_oen[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 63.280 504.000 63.880 ;
    END
  END digital_io_oen[7]
  PIN digital_io_oen[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 71.440 504.000 72.040 ;
    END
  END digital_io_oen[8]
  PIN digital_io_oen[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 79.600 504.000 80.200 ;
    END
  END digital_io_oen[9]
  PIN digital_io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 3.440 504.000 4.040 ;
    END
  END digital_io_out[0]
  PIN digital_io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 85.040 504.000 85.640 ;
    END
  END digital_io_out[10]
  PIN digital_io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 93.200 504.000 93.800 ;
    END
  END digital_io_out[11]
  PIN digital_io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 101.360 504.000 101.960 ;
    END
  END digital_io_out[12]
  PIN digital_io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 109.520 504.000 110.120 ;
    END
  END digital_io_out[13]
  PIN digital_io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 117.680 504.000 118.280 ;
    END
  END digital_io_out[14]
  PIN digital_io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 496.000 323.750 504.000 ;
    END
  END digital_io_out[15]
  PIN digital_io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 496.000 320.990 504.000 ;
    END
  END digital_io_out[16]
  PIN digital_io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 496.000 318.230 504.000 ;
    END
  END digital_io_out[17]
  PIN digital_io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 496.000 315.470 504.000 ;
    END
  END digital_io_out[18]
  PIN digital_io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 496.000 312.710 504.000 ;
    END
  END digital_io_out[19]
  PIN digital_io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 11.600 504.000 12.200 ;
    END
  END digital_io_out[1]
  PIN digital_io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 496.000 309.950 504.000 ;
    END
  END digital_io_out[20]
  PIN digital_io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 496.000 307.190 504.000 ;
    END
  END digital_io_out[21]
  PIN digital_io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 496.000 304.430 504.000 ;
    END
  END digital_io_out[22]
  PIN digital_io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 496.000 301.670 504.000 ;
    END
  END digital_io_out[23]
  PIN digital_io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 216.960 4.000 217.560 ;
    END
  END digital_io_out[24]
  PIN digital_io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 212.880 4.000 213.480 ;
    END
  END digital_io_out[25]
  PIN digital_io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 208.800 4.000 209.400 ;
    END
  END digital_io_out[26]
  PIN digital_io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 204.720 4.000 205.320 ;
    END
  END digital_io_out[27]
  PIN digital_io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 200.640 4.000 201.240 ;
    END
  END digital_io_out[28]
  PIN digital_io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 53.760 4.000 54.360 ;
    END
  END digital_io_out[29]
  PIN digital_io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 19.760 504.000 20.360 ;
    END
  END digital_io_out[2]
  PIN digital_io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 49.680 4.000 50.280 ;
    END
  END digital_io_out[30]
  PIN digital_io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 45.600 4.000 46.200 ;
    END
  END digital_io_out[31]
  PIN digital_io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 41.520 4.000 42.120 ;
    END
  END digital_io_out[32]
  PIN digital_io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 37.440 4.000 38.040 ;
    END
  END digital_io_out[33]
  PIN digital_io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 33.360 4.000 33.960 ;
    END
  END digital_io_out[34]
  PIN digital_io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 29.280 4.000 29.880 ;
    END
  END digital_io_out[35]
  PIN digital_io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 25.200 4.000 25.800 ;
    END
  END digital_io_out[36]
  PIN digital_io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 21.120 4.000 21.720 ;
    END
  END digital_io_out[37]
  PIN digital_io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 27.920 504.000 28.520 ;
    END
  END digital_io_out[3]
  PIN digital_io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 36.080 504.000 36.680 ;
    END
  END digital_io_out[4]
  PIN digital_io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 44.240 504.000 44.840 ;
    END
  END digital_io_out[5]
  PIN digital_io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 52.400 504.000 53.000 ;
    END
  END digital_io_out[6]
  PIN digital_io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 60.560 504.000 61.160 ;
    END
  END digital_io_out[7]
  PIN digital_io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 68.720 504.000 69.320 ;
    END
  END digital_io_out[8]
  PIN digital_io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 76.880 504.000 77.480 ;
    END
  END digital_io_out[9]
  PIN fuse_mhartid[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 496.000 49.590 504.000 ;
    END
  END fuse_mhartid[0]
  PIN fuse_mhartid[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 496.000 40.390 504.000 ;
    END
  END fuse_mhartid[10]
  PIN fuse_mhartid[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 496.000 39.470 504.000 ;
    END
  END fuse_mhartid[11]
  PIN fuse_mhartid[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 496.000 38.550 504.000 ;
    END
  END fuse_mhartid[12]
  PIN fuse_mhartid[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 496.000 37.630 504.000 ;
    END
  END fuse_mhartid[13]
  PIN fuse_mhartid[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 496.000 36.710 504.000 ;
    END
  END fuse_mhartid[14]
  PIN fuse_mhartid[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 496.000 35.790 504.000 ;
    END
  END fuse_mhartid[15]
  PIN fuse_mhartid[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 496.000 34.870 504.000 ;
    END
  END fuse_mhartid[16]
  PIN fuse_mhartid[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 496.000 33.950 504.000 ;
    END
  END fuse_mhartid[17]
  PIN fuse_mhartid[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 496.000 33.030 504.000 ;
    END
  END fuse_mhartid[18]
  PIN fuse_mhartid[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 496.000 32.110 504.000 ;
    END
  END fuse_mhartid[19]
  PIN fuse_mhartid[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 496.000 48.670 504.000 ;
    END
  END fuse_mhartid[1]
  PIN fuse_mhartid[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 496.000 31.190 504.000 ;
    END
  END fuse_mhartid[20]
  PIN fuse_mhartid[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 496.000 30.270 504.000 ;
    END
  END fuse_mhartid[21]
  PIN fuse_mhartid[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 496.000 29.350 504.000 ;
    END
  END fuse_mhartid[22]
  PIN fuse_mhartid[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 496.000 28.430 504.000 ;
    END
  END fuse_mhartid[23]
  PIN fuse_mhartid[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 496.000 27.510 504.000 ;
    END
  END fuse_mhartid[24]
  PIN fuse_mhartid[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 496.000 26.590 504.000 ;
    END
  END fuse_mhartid[25]
  PIN fuse_mhartid[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 496.000 25.670 504.000 ;
    END
  END fuse_mhartid[26]
  PIN fuse_mhartid[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 496.000 24.750 504.000 ;
    END
  END fuse_mhartid[27]
  PIN fuse_mhartid[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 496.000 23.830 504.000 ;
    END
  END fuse_mhartid[28]
  PIN fuse_mhartid[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 496.000 22.910 504.000 ;
    END
  END fuse_mhartid[29]
  PIN fuse_mhartid[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 496.000 47.750 504.000 ;
    END
  END fuse_mhartid[2]
  PIN fuse_mhartid[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 496.000 21.990 504.000 ;
    END
  END fuse_mhartid[30]
  PIN fuse_mhartid[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 496.000 21.070 504.000 ;
    END
  END fuse_mhartid[31]
  PIN fuse_mhartid[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 496.000 46.830 504.000 ;
    END
  END fuse_mhartid[3]
  PIN fuse_mhartid[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 496.000 45.910 504.000 ;
    END
  END fuse_mhartid[4]
  PIN fuse_mhartid[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 496.000 44.990 504.000 ;
    END
  END fuse_mhartid[5]
  PIN fuse_mhartid[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 496.000 44.070 504.000 ;
    END
  END fuse_mhartid[6]
  PIN fuse_mhartid[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 496.000 43.150 504.000 ;
    END
  END fuse_mhartid[7]
  PIN fuse_mhartid[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 496.000 42.230 504.000 ;
    END
  END fuse_mhartid[8]
  PIN fuse_mhartid[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 496.000 41.310 504.000 ;
    END
  END fuse_mhartid[9]
  PIN h_reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 496.000 1.750 504.000 ;
    END
  END h_reset_n
  PIN i2cm_clk_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 496.000 70.750 504.000 ;
    END
  END i2cm_clk_i
  PIN i2cm_clk_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 496.000 69.830 504.000 ;
    END
  END i2cm_clk_o
  PIN i2cm_clk_oen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 496.000 71.670 504.000 ;
    END
  END i2cm_clk_oen
  PIN i2cm_data_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 496.000 74.430 504.000 ;
    END
  END i2cm_data_i
  PIN i2cm_data_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 496.000 73.510 504.000 ;
    END
  END i2cm_data_o
  PIN i2cm_data_oen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 496.000 72.590 504.000 ;
    END
  END i2cm_data_oen
  PIN i2cm_intr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 496.000 79.950 504.000 ;
    END
  END i2cm_intr
  PIN irq_lines[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 496.000 16.470 504.000 ;
    END
  END irq_lines[0]
  PIN irq_lines[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 496.000 7.270 504.000 ;
    END
  END irq_lines[10]
  PIN irq_lines[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 496.000 6.350 504.000 ;
    END
  END irq_lines[11]
  PIN irq_lines[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 496.000 5.430 504.000 ;
    END
  END irq_lines[12]
  PIN irq_lines[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 496.000 4.510 504.000 ;
    END
  END irq_lines[13]
  PIN irq_lines[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 496.000 3.590 504.000 ;
    END
  END irq_lines[14]
  PIN irq_lines[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 496.000 2.670 504.000 ;
    END
  END irq_lines[15]
  PIN irq_lines[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 496.000 15.550 504.000 ;
    END
  END irq_lines[1]
  PIN irq_lines[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 496.000 14.630 504.000 ;
    END
  END irq_lines[2]
  PIN irq_lines[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 496.000 13.710 504.000 ;
    END
  END irq_lines[3]
  PIN irq_lines[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 496.000 12.790 504.000 ;
    END
  END irq_lines[4]
  PIN irq_lines[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 496.000 11.870 504.000 ;
    END
  END irq_lines[5]
  PIN irq_lines[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 496.000 10.950 504.000 ;
    END
  END irq_lines[6]
  PIN irq_lines[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 496.000 10.030 504.000 ;
    END
  END irq_lines[7]
  PIN irq_lines[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 496.000 9.110 504.000 ;
    END
  END irq_lines[8]
  PIN irq_lines[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 496.000 8.190 504.000 ;
    END
  END irq_lines[9]
  PIN mclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 496.000 0.830 504.000 ;
    END
  END mclk
  PIN pinmux_debug[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 -4.000 0.830 4.000 ;
    END
  END pinmux_debug[0]
  PIN pinmux_debug[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 -4.000 19.230 4.000 ;
    END
  END pinmux_debug[10]
  PIN pinmux_debug[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 -4.000 21.070 4.000 ;
    END
  END pinmux_debug[11]
  PIN pinmux_debug[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 -4.000 22.910 4.000 ;
    END
  END pinmux_debug[12]
  PIN pinmux_debug[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 -4.000 24.750 4.000 ;
    END
  END pinmux_debug[13]
  PIN pinmux_debug[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 -4.000 26.590 4.000 ;
    END
  END pinmux_debug[14]
  PIN pinmux_debug[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 -4.000 28.430 4.000 ;
    END
  END pinmux_debug[15]
  PIN pinmux_debug[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 -4.000 30.270 4.000 ;
    END
  END pinmux_debug[16]
  PIN pinmux_debug[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 -4.000 32.110 4.000 ;
    END
  END pinmux_debug[17]
  PIN pinmux_debug[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 -4.000 33.950 4.000 ;
    END
  END pinmux_debug[18]
  PIN pinmux_debug[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 -4.000 35.790 4.000 ;
    END
  END pinmux_debug[19]
  PIN pinmux_debug[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 -4.000 2.670 4.000 ;
    END
  END pinmux_debug[1]
  PIN pinmux_debug[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 -4.000 37.630 4.000 ;
    END
  END pinmux_debug[20]
  PIN pinmux_debug[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 -4.000 39.470 4.000 ;
    END
  END pinmux_debug[21]
  PIN pinmux_debug[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 -4.000 41.310 4.000 ;
    END
  END pinmux_debug[22]
  PIN pinmux_debug[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 -4.000 43.150 4.000 ;
    END
  END pinmux_debug[23]
  PIN pinmux_debug[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 -4.000 44.990 4.000 ;
    END
  END pinmux_debug[24]
  PIN pinmux_debug[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 -4.000 46.830 4.000 ;
    END
  END pinmux_debug[25]
  PIN pinmux_debug[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 -4.000 48.670 4.000 ;
    END
  END pinmux_debug[26]
  PIN pinmux_debug[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 -4.000 50.510 4.000 ;
    END
  END pinmux_debug[27]
  PIN pinmux_debug[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 -4.000 52.350 4.000 ;
    END
  END pinmux_debug[28]
  PIN pinmux_debug[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 -4.000 54.190 4.000 ;
    END
  END pinmux_debug[29]
  PIN pinmux_debug[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 -4.000 4.510 4.000 ;
    END
  END pinmux_debug[2]
  PIN pinmux_debug[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 -4.000 56.030 4.000 ;
    END
  END pinmux_debug[30]
  PIN pinmux_debug[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 -4.000 57.870 4.000 ;
    END
  END pinmux_debug[31]
  PIN pinmux_debug[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 -4.000 6.350 4.000 ;
    END
  END pinmux_debug[3]
  PIN pinmux_debug[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 -4.000 8.190 4.000 ;
    END
  END pinmux_debug[4]
  PIN pinmux_debug[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 -4.000 10.030 4.000 ;
    END
  END pinmux_debug[5]
  PIN pinmux_debug[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 -4.000 11.870 4.000 ;
    END
  END pinmux_debug[6]
  PIN pinmux_debug[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 -4.000 13.710 4.000 ;
    END
  END pinmux_debug[7]
  PIN pinmux_debug[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 -4.000 15.550 4.000 ;
    END
  END pinmux_debug[8]
  PIN pinmux_debug[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 -4.000 17.390 4.000 ;
    END
  END pinmux_debug[9]
  PIN pulse1m_mclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 496.000 79.030 504.000 ;
    END
  END pulse1m_mclk
  PIN reg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 496.000 272.230 504.000 ;
    END
  END reg_ack
  PIN reg_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 496.000 208.750 504.000 ;
    END
  END reg_addr[0]
  PIN reg_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 496.000 207.830 504.000 ;
    END
  END reg_addr[1]
  PIN reg_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 496.000 206.910 504.000 ;
    END
  END reg_addr[2]
  PIN reg_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 496.000 205.990 504.000 ;
    END
  END reg_addr[3]
  PIN reg_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 496.000 205.070 504.000 ;
    END
  END reg_addr[4]
  PIN reg_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 496.000 204.150 504.000 ;
    END
  END reg_addr[5]
  PIN reg_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 496.000 203.230 504.000 ;
    END
  END reg_addr[6]
  PIN reg_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 496.000 202.310 504.000 ;
    END
  END reg_addr[7]
  PIN reg_be[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 496.000 212.430 504.000 ;
    END
  END reg_be[0]
  PIN reg_be[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 496.000 211.510 504.000 ;
    END
  END reg_be[1]
  PIN reg_be[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 496.000 210.590 504.000 ;
    END
  END reg_be[2]
  PIN reg_be[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 496.000 209.670 504.000 ;
    END
  END reg_be[3]
  PIN reg_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 496.000 200.470 504.000 ;
    END
  END reg_cs
  PIN reg_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 496.000 271.310 504.000 ;
    END
  END reg_rdata[0]
  PIN reg_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 496.000 262.110 504.000 ;
    END
  END reg_rdata[10]
  PIN reg_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 496.000 261.190 504.000 ;
    END
  END reg_rdata[11]
  PIN reg_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 496.000 260.270 504.000 ;
    END
  END reg_rdata[12]
  PIN reg_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 496.000 259.350 504.000 ;
    END
  END reg_rdata[13]
  PIN reg_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 496.000 258.430 504.000 ;
    END
  END reg_rdata[14]
  PIN reg_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 496.000 257.510 504.000 ;
    END
  END reg_rdata[15]
  PIN reg_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 496.000 256.590 504.000 ;
    END
  END reg_rdata[16]
  PIN reg_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 496.000 255.670 504.000 ;
    END
  END reg_rdata[17]
  PIN reg_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 496.000 254.750 504.000 ;
    END
  END reg_rdata[18]
  PIN reg_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 496.000 253.830 504.000 ;
    END
  END reg_rdata[19]
  PIN reg_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 496.000 270.390 504.000 ;
    END
  END reg_rdata[1]
  PIN reg_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 496.000 252.910 504.000 ;
    END
  END reg_rdata[20]
  PIN reg_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 496.000 251.990 504.000 ;
    END
  END reg_rdata[21]
  PIN reg_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 496.000 251.070 504.000 ;
    END
  END reg_rdata[22]
  PIN reg_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 496.000 250.150 504.000 ;
    END
  END reg_rdata[23]
  PIN reg_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 496.000 249.230 504.000 ;
    END
  END reg_rdata[24]
  PIN reg_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 496.000 248.310 504.000 ;
    END
  END reg_rdata[25]
  PIN reg_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 496.000 247.390 504.000 ;
    END
  END reg_rdata[26]
  PIN reg_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 496.000 246.470 504.000 ;
    END
  END reg_rdata[27]
  PIN reg_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 496.000 245.550 504.000 ;
    END
  END reg_rdata[28]
  PIN reg_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 496.000 244.630 504.000 ;
    END
  END reg_rdata[29]
  PIN reg_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 496.000 269.470 504.000 ;
    END
  END reg_rdata[2]
  PIN reg_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 496.000 243.710 504.000 ;
    END
  END reg_rdata[30]
  PIN reg_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 496.000 242.790 504.000 ;
    END
  END reg_rdata[31]
  PIN reg_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 496.000 268.550 504.000 ;
    END
  END reg_rdata[3]
  PIN reg_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 496.000 267.630 504.000 ;
    END
  END reg_rdata[4]
  PIN reg_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 496.000 266.710 504.000 ;
    END
  END reg_rdata[5]
  PIN reg_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 496.000 265.790 504.000 ;
    END
  END reg_rdata[6]
  PIN reg_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 496.000 264.870 504.000 ;
    END
  END reg_rdata[7]
  PIN reg_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 496.000 263.950 504.000 ;
    END
  END reg_rdata[8]
  PIN reg_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 496.000 263.030 504.000 ;
    END
  END reg_rdata[9]
  PIN reg_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 496.000 241.870 504.000 ;
    END
  END reg_wdata[0]
  PIN reg_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 496.000 232.670 504.000 ;
    END
  END reg_wdata[10]
  PIN reg_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 496.000 231.750 504.000 ;
    END
  END reg_wdata[11]
  PIN reg_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 496.000 230.830 504.000 ;
    END
  END reg_wdata[12]
  PIN reg_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 496.000 229.910 504.000 ;
    END
  END reg_wdata[13]
  PIN reg_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 496.000 228.990 504.000 ;
    END
  END reg_wdata[14]
  PIN reg_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 496.000 228.070 504.000 ;
    END
  END reg_wdata[15]
  PIN reg_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 496.000 227.150 504.000 ;
    END
  END reg_wdata[16]
  PIN reg_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 496.000 226.230 504.000 ;
    END
  END reg_wdata[17]
  PIN reg_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 496.000 225.310 504.000 ;
    END
  END reg_wdata[18]
  PIN reg_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 496.000 224.390 504.000 ;
    END
  END reg_wdata[19]
  PIN reg_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 496.000 240.950 504.000 ;
    END
  END reg_wdata[1]
  PIN reg_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 496.000 223.470 504.000 ;
    END
  END reg_wdata[20]
  PIN reg_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 496.000 222.550 504.000 ;
    END
  END reg_wdata[21]
  PIN reg_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 496.000 221.630 504.000 ;
    END
  END reg_wdata[22]
  PIN reg_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 496.000 220.710 504.000 ;
    END
  END reg_wdata[23]
  PIN reg_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 496.000 219.790 504.000 ;
    END
  END reg_wdata[24]
  PIN reg_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 496.000 218.870 504.000 ;
    END
  END reg_wdata[25]
  PIN reg_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 496.000 217.950 504.000 ;
    END
  END reg_wdata[26]
  PIN reg_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 496.000 217.030 504.000 ;
    END
  END reg_wdata[27]
  PIN reg_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 496.000 216.110 504.000 ;
    END
  END reg_wdata[28]
  PIN reg_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 496.000 215.190 504.000 ;
    END
  END reg_wdata[29]
  PIN reg_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 496.000 240.030 504.000 ;
    END
  END reg_wdata[2]
  PIN reg_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 496.000 214.270 504.000 ;
    END
  END reg_wdata[30]
  PIN reg_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 496.000 213.350 504.000 ;
    END
  END reg_wdata[31]
  PIN reg_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 496.000 239.110 504.000 ;
    END
  END reg_wdata[3]
  PIN reg_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 496.000 238.190 504.000 ;
    END
  END reg_wdata[4]
  PIN reg_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 496.000 237.270 504.000 ;
    END
  END reg_wdata[5]
  PIN reg_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 496.000 236.350 504.000 ;
    END
  END reg_wdata[6]
  PIN reg_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 496.000 235.430 504.000 ;
    END
  END reg_wdata[7]
  PIN reg_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 496.000 234.510 504.000 ;
    END
  END reg_wdata[8]
  PIN reg_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 496.000 233.590 504.000 ;
    END
  END reg_wdata[9]
  PIN reg_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 496.000 201.390 504.000 ;
    END
  END reg_wr
  PIN sflash_di[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 14.320 4.000 14.920 ;
    END
  END sflash_di[0]
  PIN sflash_di[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 15.680 4.000 16.280 ;
    END
  END sflash_di[1]
  PIN sflash_di[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 17.040 4.000 17.640 ;
    END
  END sflash_di[2]
  PIN sflash_di[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 18.400 4.000 19.000 ;
    END
  END sflash_di[3]
  PIN sflash_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 8.880 4.000 9.480 ;
    END
  END sflash_do[0]
  PIN sflash_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 10.240 4.000 10.840 ;
    END
  END sflash_do[1]
  PIN sflash_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 11.600 4.000 12.200 ;
    END
  END sflash_do[2]
  PIN sflash_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 12.960 4.000 13.560 ;
    END
  END sflash_do[3]
  PIN sflash_oen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 0.720 4.000 1.320 ;
    END
  END sflash_oen[0]
  PIN sflash_oen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2.080 4.000 2.680 ;
    END
  END sflash_oen[1]
  PIN sflash_oen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 3.440 4.000 4.040 ;
    END
  END sflash_oen[2]
  PIN sflash_oen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 4.800 4.000 5.400 ;
    END
  END sflash_oen[3]
  PIN sflash_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 7.520 4.000 8.120 ;
    END
  END sflash_sck
  PIN sflash_ss
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 6.160 4.000 6.760 ;
    END
  END sflash_ss
  PIN soft_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 496.000 20.150 504.000 ;
    END
  END soft_irq
  PIN spim_miso
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 496.000 77.190 504.000 ;
    END
  END spim_miso
  PIN spim_mosi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 496.000 78.110 504.000 ;
    END
  END spim_mosi
  PIN spim_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 496.000 75.350 504.000 ;
    END
  END spim_sck
  PIN spim_ss
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 496.000 76.270 504.000 ;
    END
  END spim_ss
  PIN ssram_di[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 496.000 62.470 504.000 ;
    END
  END ssram_di[0]
  PIN ssram_di[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 496.000 61.550 504.000 ;
    END
  END ssram_di[1]
  PIN ssram_di[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 496.000 60.630 504.000 ;
    END
  END ssram_di[2]
  PIN ssram_di[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 496.000 59.710 504.000 ;
    END
  END ssram_di[3]
  PIN ssram_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 496.000 58.790 504.000 ;
    END
  END ssram_do[0]
  PIN ssram_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 496.000 57.870 504.000 ;
    END
  END ssram_do[1]
  PIN ssram_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 496.000 56.950 504.000 ;
    END
  END ssram_do[2]
  PIN ssram_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 496.000 56.030 504.000 ;
    END
  END ssram_do[3]
  PIN ssram_oen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 496.000 55.110 504.000 ;
    END
  END ssram_oen[0]
  PIN ssram_oen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 496.000 54.190 504.000 ;
    END
  END ssram_oen[1]
  PIN ssram_oen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 496.000 53.270 504.000 ;
    END
  END ssram_oen[2]
  PIN ssram_oen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 496.000 52.350 504.000 ;
    END
  END ssram_oen[3]
  PIN ssram_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 496.000 50.510 504.000 ;
    END
  END ssram_sck
  PIN ssram_ss
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 496.000 51.430 504.000 ;
    END
  END ssram_ss
  PIN uart_rxd
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 496.000 68.910 504.000 ;
    END
  END uart_rxd
  PIN uart_txd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 496.000 67.990 504.000 ;
    END
  END uart_txd
  PIN usb_dn_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 496.000 67.070 504.000 ;
    END
  END usb_dn_i
  PIN usb_dn_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 496.000 64.310 504.000 ;
    END
  END usb_dn_o
  PIN usb_dp_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 496.000 66.150 504.000 ;
    END
  END usb_dp_i
  PIN usb_dp_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 496.000 63.390 504.000 ;
    END
  END usb_dp_o
  PIN usb_intr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 496.000 80.870 504.000 ;
    END
  END usb_intr
  PIN usb_oen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 496.000 65.230 504.000 ;
    END
  END usb_oen
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 496.000 19.230 504.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 496.000 18.310 504.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 496.000 17.390 504.000 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.340 10.640 24.340 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.340 10.640 124.340 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 219.340 10.640 224.340 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 319.340 10.640 324.340 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 419.340 10.640 424.340 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 69.340 10.640 74.340 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 169.340 10.640 174.340 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 269.340 10.640 274.340 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 369.340 10.640 374.340 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 469.340 10.640 474.340 487.120 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.815 489.855 ;
      LAYER met1 ;
        RECT 0.530 2.420 494.875 491.260 ;
      LAYER met2 ;
        RECT 1.110 495.720 1.190 496.000 ;
        RECT 2.030 495.720 2.110 496.000 ;
        RECT 2.950 495.720 3.030 496.000 ;
        RECT 3.870 495.720 3.950 496.000 ;
        RECT 4.790 495.720 4.870 496.000 ;
        RECT 5.710 495.720 5.790 496.000 ;
        RECT 6.630 495.720 6.710 496.000 ;
        RECT 7.550 495.720 7.630 496.000 ;
        RECT 8.470 495.720 8.550 496.000 ;
        RECT 9.390 495.720 9.470 496.000 ;
        RECT 10.310 495.720 10.390 496.000 ;
        RECT 11.230 495.720 11.310 496.000 ;
        RECT 12.150 495.720 12.230 496.000 ;
        RECT 13.070 495.720 13.150 496.000 ;
        RECT 13.990 495.720 14.070 496.000 ;
        RECT 14.910 495.720 14.990 496.000 ;
        RECT 15.830 495.720 15.910 496.000 ;
        RECT 16.750 495.720 16.830 496.000 ;
        RECT 17.670 495.720 17.750 496.000 ;
        RECT 18.590 495.720 18.670 496.000 ;
        RECT 19.510 495.720 19.590 496.000 ;
        RECT 20.430 495.720 20.510 496.000 ;
        RECT 21.350 495.720 21.430 496.000 ;
        RECT 22.270 495.720 22.350 496.000 ;
        RECT 23.190 495.720 23.270 496.000 ;
        RECT 24.110 495.720 24.190 496.000 ;
        RECT 25.030 495.720 25.110 496.000 ;
        RECT 25.950 495.720 26.030 496.000 ;
        RECT 26.870 495.720 26.950 496.000 ;
        RECT 27.790 495.720 27.870 496.000 ;
        RECT 28.710 495.720 28.790 496.000 ;
        RECT 29.630 495.720 29.710 496.000 ;
        RECT 30.550 495.720 30.630 496.000 ;
        RECT 31.470 495.720 31.550 496.000 ;
        RECT 32.390 495.720 32.470 496.000 ;
        RECT 33.310 495.720 33.390 496.000 ;
        RECT 34.230 495.720 34.310 496.000 ;
        RECT 35.150 495.720 35.230 496.000 ;
        RECT 36.070 495.720 36.150 496.000 ;
        RECT 36.990 495.720 37.070 496.000 ;
        RECT 37.910 495.720 37.990 496.000 ;
        RECT 38.830 495.720 38.910 496.000 ;
        RECT 39.750 495.720 39.830 496.000 ;
        RECT 40.670 495.720 40.750 496.000 ;
        RECT 41.590 495.720 41.670 496.000 ;
        RECT 42.510 495.720 42.590 496.000 ;
        RECT 43.430 495.720 43.510 496.000 ;
        RECT 44.350 495.720 44.430 496.000 ;
        RECT 45.270 495.720 45.350 496.000 ;
        RECT 46.190 495.720 46.270 496.000 ;
        RECT 47.110 495.720 47.190 496.000 ;
        RECT 48.030 495.720 48.110 496.000 ;
        RECT 48.950 495.720 49.030 496.000 ;
        RECT 49.870 495.720 49.950 496.000 ;
        RECT 50.790 495.720 50.870 496.000 ;
        RECT 51.710 495.720 51.790 496.000 ;
        RECT 52.630 495.720 52.710 496.000 ;
        RECT 53.550 495.720 53.630 496.000 ;
        RECT 54.470 495.720 54.550 496.000 ;
        RECT 55.390 495.720 55.470 496.000 ;
        RECT 56.310 495.720 56.390 496.000 ;
        RECT 57.230 495.720 57.310 496.000 ;
        RECT 58.150 495.720 58.230 496.000 ;
        RECT 59.070 495.720 59.150 496.000 ;
        RECT 59.990 495.720 60.070 496.000 ;
        RECT 60.910 495.720 60.990 496.000 ;
        RECT 61.830 495.720 61.910 496.000 ;
        RECT 62.750 495.720 62.830 496.000 ;
        RECT 63.670 495.720 63.750 496.000 ;
        RECT 64.590 495.720 64.670 496.000 ;
        RECT 65.510 495.720 65.590 496.000 ;
        RECT 66.430 495.720 66.510 496.000 ;
        RECT 67.350 495.720 67.430 496.000 ;
        RECT 68.270 495.720 68.350 496.000 ;
        RECT 69.190 495.720 69.270 496.000 ;
        RECT 70.110 495.720 70.190 496.000 ;
        RECT 71.030 495.720 71.110 496.000 ;
        RECT 71.950 495.720 72.030 496.000 ;
        RECT 72.870 495.720 72.950 496.000 ;
        RECT 73.790 495.720 73.870 496.000 ;
        RECT 74.710 495.720 74.790 496.000 ;
        RECT 75.630 495.720 75.710 496.000 ;
        RECT 76.550 495.720 76.630 496.000 ;
        RECT 77.470 495.720 77.550 496.000 ;
        RECT 78.390 495.720 78.470 496.000 ;
        RECT 79.310 495.720 79.390 496.000 ;
        RECT 80.230 495.720 80.310 496.000 ;
        RECT 81.150 495.720 199.910 496.000 ;
        RECT 200.750 495.720 200.830 496.000 ;
        RECT 201.670 495.720 201.750 496.000 ;
        RECT 202.590 495.720 202.670 496.000 ;
        RECT 203.510 495.720 203.590 496.000 ;
        RECT 204.430 495.720 204.510 496.000 ;
        RECT 205.350 495.720 205.430 496.000 ;
        RECT 206.270 495.720 206.350 496.000 ;
        RECT 207.190 495.720 207.270 496.000 ;
        RECT 208.110 495.720 208.190 496.000 ;
        RECT 209.030 495.720 209.110 496.000 ;
        RECT 209.950 495.720 210.030 496.000 ;
        RECT 210.870 495.720 210.950 496.000 ;
        RECT 211.790 495.720 211.870 496.000 ;
        RECT 212.710 495.720 212.790 496.000 ;
        RECT 213.630 495.720 213.710 496.000 ;
        RECT 214.550 495.720 214.630 496.000 ;
        RECT 215.470 495.720 215.550 496.000 ;
        RECT 216.390 495.720 216.470 496.000 ;
        RECT 217.310 495.720 217.390 496.000 ;
        RECT 218.230 495.720 218.310 496.000 ;
        RECT 219.150 495.720 219.230 496.000 ;
        RECT 220.070 495.720 220.150 496.000 ;
        RECT 220.990 495.720 221.070 496.000 ;
        RECT 221.910 495.720 221.990 496.000 ;
        RECT 222.830 495.720 222.910 496.000 ;
        RECT 223.750 495.720 223.830 496.000 ;
        RECT 224.670 495.720 224.750 496.000 ;
        RECT 225.590 495.720 225.670 496.000 ;
        RECT 226.510 495.720 226.590 496.000 ;
        RECT 227.430 495.720 227.510 496.000 ;
        RECT 228.350 495.720 228.430 496.000 ;
        RECT 229.270 495.720 229.350 496.000 ;
        RECT 230.190 495.720 230.270 496.000 ;
        RECT 231.110 495.720 231.190 496.000 ;
        RECT 232.030 495.720 232.110 496.000 ;
        RECT 232.950 495.720 233.030 496.000 ;
        RECT 233.870 495.720 233.950 496.000 ;
        RECT 234.790 495.720 234.870 496.000 ;
        RECT 235.710 495.720 235.790 496.000 ;
        RECT 236.630 495.720 236.710 496.000 ;
        RECT 237.550 495.720 237.630 496.000 ;
        RECT 238.470 495.720 238.550 496.000 ;
        RECT 239.390 495.720 239.470 496.000 ;
        RECT 240.310 495.720 240.390 496.000 ;
        RECT 241.230 495.720 241.310 496.000 ;
        RECT 242.150 495.720 242.230 496.000 ;
        RECT 243.070 495.720 243.150 496.000 ;
        RECT 243.990 495.720 244.070 496.000 ;
        RECT 244.910 495.720 244.990 496.000 ;
        RECT 245.830 495.720 245.910 496.000 ;
        RECT 246.750 495.720 246.830 496.000 ;
        RECT 247.670 495.720 247.750 496.000 ;
        RECT 248.590 495.720 248.670 496.000 ;
        RECT 249.510 495.720 249.590 496.000 ;
        RECT 250.430 495.720 250.510 496.000 ;
        RECT 251.350 495.720 251.430 496.000 ;
        RECT 252.270 495.720 252.350 496.000 ;
        RECT 253.190 495.720 253.270 496.000 ;
        RECT 254.110 495.720 254.190 496.000 ;
        RECT 255.030 495.720 255.110 496.000 ;
        RECT 255.950 495.720 256.030 496.000 ;
        RECT 256.870 495.720 256.950 496.000 ;
        RECT 257.790 495.720 257.870 496.000 ;
        RECT 258.710 495.720 258.790 496.000 ;
        RECT 259.630 495.720 259.710 496.000 ;
        RECT 260.550 495.720 260.630 496.000 ;
        RECT 261.470 495.720 261.550 496.000 ;
        RECT 262.390 495.720 262.470 496.000 ;
        RECT 263.310 495.720 263.390 496.000 ;
        RECT 264.230 495.720 264.310 496.000 ;
        RECT 265.150 495.720 265.230 496.000 ;
        RECT 266.070 495.720 266.150 496.000 ;
        RECT 266.990 495.720 267.070 496.000 ;
        RECT 267.910 495.720 267.990 496.000 ;
        RECT 268.830 495.720 268.910 496.000 ;
        RECT 269.750 495.720 269.830 496.000 ;
        RECT 270.670 495.720 270.750 496.000 ;
        RECT 271.590 495.720 271.670 496.000 ;
        RECT 272.510 495.720 300.190 496.000 ;
        RECT 301.030 495.720 301.110 496.000 ;
        RECT 301.950 495.720 302.030 496.000 ;
        RECT 302.870 495.720 302.950 496.000 ;
        RECT 303.790 495.720 303.870 496.000 ;
        RECT 304.710 495.720 304.790 496.000 ;
        RECT 305.630 495.720 305.710 496.000 ;
        RECT 306.550 495.720 306.630 496.000 ;
        RECT 307.470 495.720 307.550 496.000 ;
        RECT 308.390 495.720 308.470 496.000 ;
        RECT 309.310 495.720 309.390 496.000 ;
        RECT 310.230 495.720 310.310 496.000 ;
        RECT 311.150 495.720 311.230 496.000 ;
        RECT 312.070 495.720 312.150 496.000 ;
        RECT 312.990 495.720 313.070 496.000 ;
        RECT 313.910 495.720 313.990 496.000 ;
        RECT 314.830 495.720 314.910 496.000 ;
        RECT 315.750 495.720 315.830 496.000 ;
        RECT 316.670 495.720 316.750 496.000 ;
        RECT 317.590 495.720 317.670 496.000 ;
        RECT 318.510 495.720 318.590 496.000 ;
        RECT 319.430 495.720 319.510 496.000 ;
        RECT 320.350 495.720 320.430 496.000 ;
        RECT 321.270 495.720 321.350 496.000 ;
        RECT 322.190 495.720 322.270 496.000 ;
        RECT 323.110 495.720 323.190 496.000 ;
        RECT 324.030 495.720 324.110 496.000 ;
        RECT 324.950 495.720 490.730 496.000 ;
        RECT 0.560 4.280 490.730 495.720 ;
        RECT 1.110 0.835 2.110 4.280 ;
        RECT 2.950 0.835 3.950 4.280 ;
        RECT 4.790 0.835 5.790 4.280 ;
        RECT 6.630 0.835 7.630 4.280 ;
        RECT 8.470 0.835 9.470 4.280 ;
        RECT 10.310 0.835 11.310 4.280 ;
        RECT 12.150 0.835 13.150 4.280 ;
        RECT 13.990 0.835 14.990 4.280 ;
        RECT 15.830 0.835 16.830 4.280 ;
        RECT 17.670 0.835 18.670 4.280 ;
        RECT 19.510 0.835 20.510 4.280 ;
        RECT 21.350 0.835 22.350 4.280 ;
        RECT 23.190 0.835 24.190 4.280 ;
        RECT 25.030 0.835 26.030 4.280 ;
        RECT 26.870 0.835 27.870 4.280 ;
        RECT 28.710 0.835 29.710 4.280 ;
        RECT 30.550 0.835 31.550 4.280 ;
        RECT 32.390 0.835 33.390 4.280 ;
        RECT 34.230 0.835 35.230 4.280 ;
        RECT 36.070 0.835 37.070 4.280 ;
        RECT 37.910 0.835 38.910 4.280 ;
        RECT 39.750 0.835 40.750 4.280 ;
        RECT 41.590 0.835 42.590 4.280 ;
        RECT 43.430 0.835 44.430 4.280 ;
        RECT 45.270 0.835 46.270 4.280 ;
        RECT 47.110 0.835 48.110 4.280 ;
        RECT 48.950 0.835 49.950 4.280 ;
        RECT 50.790 0.835 51.790 4.280 ;
        RECT 52.630 0.835 53.630 4.280 ;
        RECT 54.470 0.835 55.470 4.280 ;
        RECT 56.310 0.835 57.310 4.280 ;
        RECT 58.150 0.835 490.730 4.280 ;
      LAYER met3 ;
        RECT 2.365 219.320 496.000 488.065 ;
        RECT 4.400 200.240 496.000 219.320 ;
        RECT 2.365 121.400 496.000 200.240 ;
        RECT 2.365 120.000 495.600 121.400 ;
        RECT 2.365 118.680 496.000 120.000 ;
        RECT 2.365 117.280 495.600 118.680 ;
        RECT 2.365 115.960 496.000 117.280 ;
        RECT 2.365 114.560 495.600 115.960 ;
        RECT 2.365 113.240 496.000 114.560 ;
        RECT 2.365 111.840 495.600 113.240 ;
        RECT 2.365 110.520 496.000 111.840 ;
        RECT 2.365 109.120 495.600 110.520 ;
        RECT 2.365 107.800 496.000 109.120 ;
        RECT 2.365 106.400 495.600 107.800 ;
        RECT 2.365 105.080 496.000 106.400 ;
        RECT 2.365 103.680 495.600 105.080 ;
        RECT 2.365 102.360 496.000 103.680 ;
        RECT 2.365 100.960 495.600 102.360 ;
        RECT 2.365 99.640 496.000 100.960 ;
        RECT 2.365 98.240 495.600 99.640 ;
        RECT 2.365 96.920 496.000 98.240 ;
        RECT 2.365 95.520 495.600 96.920 ;
        RECT 2.365 94.200 496.000 95.520 ;
        RECT 2.365 92.800 495.600 94.200 ;
        RECT 2.365 91.480 496.000 92.800 ;
        RECT 2.365 90.080 495.600 91.480 ;
        RECT 2.365 88.760 496.000 90.080 ;
        RECT 2.365 87.360 495.600 88.760 ;
        RECT 2.365 86.040 496.000 87.360 ;
        RECT 2.365 84.640 495.600 86.040 ;
        RECT 2.365 83.320 496.000 84.640 ;
        RECT 2.365 81.920 495.600 83.320 ;
        RECT 2.365 80.600 496.000 81.920 ;
        RECT 2.365 79.200 495.600 80.600 ;
        RECT 2.365 77.880 496.000 79.200 ;
        RECT 2.365 76.480 495.600 77.880 ;
        RECT 2.365 75.160 496.000 76.480 ;
        RECT 2.365 73.760 495.600 75.160 ;
        RECT 2.365 72.440 496.000 73.760 ;
        RECT 2.365 71.040 495.600 72.440 ;
        RECT 2.365 69.720 496.000 71.040 ;
        RECT 2.365 68.320 495.600 69.720 ;
        RECT 2.365 67.000 496.000 68.320 ;
        RECT 2.365 65.600 495.600 67.000 ;
        RECT 2.365 64.280 496.000 65.600 ;
        RECT 2.365 62.880 495.600 64.280 ;
        RECT 2.365 61.560 496.000 62.880 ;
        RECT 2.365 60.160 495.600 61.560 ;
        RECT 2.365 58.840 496.000 60.160 ;
        RECT 2.365 57.480 495.600 58.840 ;
        RECT 4.400 57.440 495.600 57.480 ;
        RECT 4.400 56.120 496.000 57.440 ;
        RECT 4.400 54.720 495.600 56.120 ;
        RECT 4.400 53.400 496.000 54.720 ;
        RECT 4.400 52.000 495.600 53.400 ;
        RECT 4.400 50.680 496.000 52.000 ;
        RECT 4.400 49.280 495.600 50.680 ;
        RECT 4.400 47.960 496.000 49.280 ;
        RECT 4.400 46.560 495.600 47.960 ;
        RECT 4.400 45.240 496.000 46.560 ;
        RECT 4.400 43.840 495.600 45.240 ;
        RECT 4.400 42.520 496.000 43.840 ;
        RECT 4.400 41.120 495.600 42.520 ;
        RECT 4.400 39.800 496.000 41.120 ;
        RECT 4.400 38.400 495.600 39.800 ;
        RECT 4.400 37.080 496.000 38.400 ;
        RECT 4.400 35.680 495.600 37.080 ;
        RECT 4.400 34.360 496.000 35.680 ;
        RECT 4.400 32.960 495.600 34.360 ;
        RECT 4.400 31.640 496.000 32.960 ;
        RECT 4.400 30.240 495.600 31.640 ;
        RECT 4.400 28.920 496.000 30.240 ;
        RECT 4.400 27.520 495.600 28.920 ;
        RECT 4.400 26.200 496.000 27.520 ;
        RECT 4.400 24.800 495.600 26.200 ;
        RECT 4.400 23.480 496.000 24.800 ;
        RECT 4.400 22.080 495.600 23.480 ;
        RECT 4.400 20.760 496.000 22.080 ;
        RECT 4.400 19.360 495.600 20.760 ;
        RECT 4.400 18.040 496.000 19.360 ;
        RECT 4.400 16.640 495.600 18.040 ;
        RECT 4.400 15.320 496.000 16.640 ;
        RECT 4.400 13.920 495.600 15.320 ;
        RECT 4.400 12.600 496.000 13.920 ;
        RECT 4.400 11.200 495.600 12.600 ;
        RECT 4.400 9.880 496.000 11.200 ;
        RECT 4.400 8.480 495.600 9.880 ;
        RECT 4.400 7.160 496.000 8.480 ;
        RECT 4.400 5.760 495.600 7.160 ;
        RECT 4.400 4.440 496.000 5.760 ;
        RECT 4.400 3.040 495.600 4.440 ;
        RECT 4.400 1.720 496.000 3.040 ;
        RECT 4.400 0.855 495.600 1.720 ;
      LAYER met4 ;
        RECT 51.815 39.615 68.940 484.665 ;
        RECT 74.740 39.615 118.940 484.665 ;
        RECT 124.740 39.615 168.940 484.665 ;
        RECT 174.740 39.615 218.940 484.665 ;
        RECT 224.740 39.615 268.940 484.665 ;
        RECT 274.740 39.615 318.940 484.665 ;
        RECT 324.740 39.615 368.940 484.665 ;
        RECT 374.740 39.615 418.940 484.665 ;
        RECT 424.740 39.615 468.940 484.665 ;
        RECT 474.740 39.615 475.345 484.665 ;
  END
END pinmux
MACRO wb_interconnect
  CLASS BLOCK ;
  FOREIGN wb_interconnect ;
  ORIGIN 0.000 0.000 ;
  SIZE 2200.000 BY 150.000 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2196.000 0.720 2204.000 1.320 ;
    END
  END clk_i
  PIN m0_wbd_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 -4.000 94.670 4.000 ;
    END
  END m0_wbd_ack_o
  PIN m0_wbd_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 -4.000 31.190 4.000 ;
    END
  END m0_wbd_adr_i[0]
  PIN m0_wbd_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 -4.000 21.990 4.000 ;
    END
  END m0_wbd_adr_i[10]
  PIN m0_wbd_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 -4.000 21.070 4.000 ;
    END
  END m0_wbd_adr_i[11]
  PIN m0_wbd_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 -4.000 20.150 4.000 ;
    END
  END m0_wbd_adr_i[12]
  PIN m0_wbd_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 -4.000 19.230 4.000 ;
    END
  END m0_wbd_adr_i[13]
  PIN m0_wbd_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 -4.000 18.310 4.000 ;
    END
  END m0_wbd_adr_i[14]
  PIN m0_wbd_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 -4.000 17.390 4.000 ;
    END
  END m0_wbd_adr_i[15]
  PIN m0_wbd_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 -4.000 16.470 4.000 ;
    END
  END m0_wbd_adr_i[16]
  PIN m0_wbd_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 -4.000 15.550 4.000 ;
    END
  END m0_wbd_adr_i[17]
  PIN m0_wbd_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 -4.000 14.630 4.000 ;
    END
  END m0_wbd_adr_i[18]
  PIN m0_wbd_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 -4.000 13.710 4.000 ;
    END
  END m0_wbd_adr_i[19]
  PIN m0_wbd_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 -4.000 30.270 4.000 ;
    END
  END m0_wbd_adr_i[1]
  PIN m0_wbd_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 -4.000 12.790 4.000 ;
    END
  END m0_wbd_adr_i[20]
  PIN m0_wbd_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 -4.000 11.870 4.000 ;
    END
  END m0_wbd_adr_i[21]
  PIN m0_wbd_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 -4.000 10.950 4.000 ;
    END
  END m0_wbd_adr_i[22]
  PIN m0_wbd_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 -4.000 10.030 4.000 ;
    END
  END m0_wbd_adr_i[23]
  PIN m0_wbd_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 -4.000 9.110 4.000 ;
    END
  END m0_wbd_adr_i[24]
  PIN m0_wbd_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 -4.000 8.190 4.000 ;
    END
  END m0_wbd_adr_i[25]
  PIN m0_wbd_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 -4.000 7.270 4.000 ;
    END
  END m0_wbd_adr_i[26]
  PIN m0_wbd_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 -4.000 6.350 4.000 ;
    END
  END m0_wbd_adr_i[27]
  PIN m0_wbd_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 -4.000 5.430 4.000 ;
    END
  END m0_wbd_adr_i[28]
  PIN m0_wbd_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 -4.000 4.510 4.000 ;
    END
  END m0_wbd_adr_i[29]
  PIN m0_wbd_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 -4.000 29.350 4.000 ;
    END
  END m0_wbd_adr_i[2]
  PIN m0_wbd_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 -4.000 3.590 4.000 ;
    END
  END m0_wbd_adr_i[30]
  PIN m0_wbd_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 -4.000 2.670 4.000 ;
    END
  END m0_wbd_adr_i[31]
  PIN m0_wbd_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 -4.000 28.430 4.000 ;
    END
  END m0_wbd_adr_i[3]
  PIN m0_wbd_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 -4.000 27.510 4.000 ;
    END
  END m0_wbd_adr_i[4]
  PIN m0_wbd_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 -4.000 26.590 4.000 ;
    END
  END m0_wbd_adr_i[5]
  PIN m0_wbd_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 -4.000 25.670 4.000 ;
    END
  END m0_wbd_adr_i[6]
  PIN m0_wbd_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 -4.000 24.750 4.000 ;
    END
  END m0_wbd_adr_i[7]
  PIN m0_wbd_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 -4.000 23.830 4.000 ;
    END
  END m0_wbd_adr_i[8]
  PIN m0_wbd_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 -4.000 22.910 4.000 ;
    END
  END m0_wbd_adr_i[9]
  PIN m0_wbd_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 -4.000 96.510 4.000 ;
    END
  END m0_wbd_cyc_i
  PIN m0_wbd_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 -4.000 64.310 4.000 ;
    END
  END m0_wbd_dat_i[0]
  PIN m0_wbd_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 -4.000 55.110 4.000 ;
    END
  END m0_wbd_dat_i[10]
  PIN m0_wbd_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 -4.000 54.190 4.000 ;
    END
  END m0_wbd_dat_i[11]
  PIN m0_wbd_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 -4.000 53.270 4.000 ;
    END
  END m0_wbd_dat_i[12]
  PIN m0_wbd_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 -4.000 52.350 4.000 ;
    END
  END m0_wbd_dat_i[13]
  PIN m0_wbd_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 -4.000 51.430 4.000 ;
    END
  END m0_wbd_dat_i[14]
  PIN m0_wbd_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 -4.000 50.510 4.000 ;
    END
  END m0_wbd_dat_i[15]
  PIN m0_wbd_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 -4.000 49.590 4.000 ;
    END
  END m0_wbd_dat_i[16]
  PIN m0_wbd_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 -4.000 48.670 4.000 ;
    END
  END m0_wbd_dat_i[17]
  PIN m0_wbd_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 -4.000 47.750 4.000 ;
    END
  END m0_wbd_dat_i[18]
  PIN m0_wbd_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 -4.000 46.830 4.000 ;
    END
  END m0_wbd_dat_i[19]
  PIN m0_wbd_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 -4.000 63.390 4.000 ;
    END
  END m0_wbd_dat_i[1]
  PIN m0_wbd_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 -4.000 45.910 4.000 ;
    END
  END m0_wbd_dat_i[20]
  PIN m0_wbd_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 -4.000 44.990 4.000 ;
    END
  END m0_wbd_dat_i[21]
  PIN m0_wbd_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 -4.000 44.070 4.000 ;
    END
  END m0_wbd_dat_i[22]
  PIN m0_wbd_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 -4.000 43.150 4.000 ;
    END
  END m0_wbd_dat_i[23]
  PIN m0_wbd_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 -4.000 42.230 4.000 ;
    END
  END m0_wbd_dat_i[24]
  PIN m0_wbd_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 -4.000 41.310 4.000 ;
    END
  END m0_wbd_dat_i[25]
  PIN m0_wbd_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 -4.000 40.390 4.000 ;
    END
  END m0_wbd_dat_i[26]
  PIN m0_wbd_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 -4.000 39.470 4.000 ;
    END
  END m0_wbd_dat_i[27]
  PIN m0_wbd_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 -4.000 38.550 4.000 ;
    END
  END m0_wbd_dat_i[28]
  PIN m0_wbd_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 -4.000 37.630 4.000 ;
    END
  END m0_wbd_dat_i[29]
  PIN m0_wbd_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 -4.000 62.470 4.000 ;
    END
  END m0_wbd_dat_i[2]
  PIN m0_wbd_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 -4.000 36.710 4.000 ;
    END
  END m0_wbd_dat_i[30]
  PIN m0_wbd_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 -4.000 35.790 4.000 ;
    END
  END m0_wbd_dat_i[31]
  PIN m0_wbd_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 -4.000 61.550 4.000 ;
    END
  END m0_wbd_dat_i[3]
  PIN m0_wbd_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 -4.000 60.630 4.000 ;
    END
  END m0_wbd_dat_i[4]
  PIN m0_wbd_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 -4.000 59.710 4.000 ;
    END
  END m0_wbd_dat_i[5]
  PIN m0_wbd_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 -4.000 58.790 4.000 ;
    END
  END m0_wbd_dat_i[6]
  PIN m0_wbd_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 -4.000 57.870 4.000 ;
    END
  END m0_wbd_dat_i[7]
  PIN m0_wbd_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 -4.000 56.950 4.000 ;
    END
  END m0_wbd_dat_i[8]
  PIN m0_wbd_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 -4.000 56.030 4.000 ;
    END
  END m0_wbd_dat_i[9]
  PIN m0_wbd_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 -4.000 93.750 4.000 ;
    END
  END m0_wbd_dat_o[0]
  PIN m0_wbd_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 -4.000 84.550 4.000 ;
    END
  END m0_wbd_dat_o[10]
  PIN m0_wbd_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 -4.000 83.630 4.000 ;
    END
  END m0_wbd_dat_o[11]
  PIN m0_wbd_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 -4.000 82.710 4.000 ;
    END
  END m0_wbd_dat_o[12]
  PIN m0_wbd_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 -4.000 81.790 4.000 ;
    END
  END m0_wbd_dat_o[13]
  PIN m0_wbd_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 -4.000 80.870 4.000 ;
    END
  END m0_wbd_dat_o[14]
  PIN m0_wbd_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 -4.000 79.950 4.000 ;
    END
  END m0_wbd_dat_o[15]
  PIN m0_wbd_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 -4.000 79.030 4.000 ;
    END
  END m0_wbd_dat_o[16]
  PIN m0_wbd_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 -4.000 78.110 4.000 ;
    END
  END m0_wbd_dat_o[17]
  PIN m0_wbd_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 -4.000 77.190 4.000 ;
    END
  END m0_wbd_dat_o[18]
  PIN m0_wbd_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 -4.000 76.270 4.000 ;
    END
  END m0_wbd_dat_o[19]
  PIN m0_wbd_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 -4.000 92.830 4.000 ;
    END
  END m0_wbd_dat_o[1]
  PIN m0_wbd_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 -4.000 75.350 4.000 ;
    END
  END m0_wbd_dat_o[20]
  PIN m0_wbd_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 -4.000 74.430 4.000 ;
    END
  END m0_wbd_dat_o[21]
  PIN m0_wbd_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 -4.000 73.510 4.000 ;
    END
  END m0_wbd_dat_o[22]
  PIN m0_wbd_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 -4.000 72.590 4.000 ;
    END
  END m0_wbd_dat_o[23]
  PIN m0_wbd_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 -4.000 71.670 4.000 ;
    END
  END m0_wbd_dat_o[24]
  PIN m0_wbd_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 -4.000 70.750 4.000 ;
    END
  END m0_wbd_dat_o[25]
  PIN m0_wbd_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 -4.000 69.830 4.000 ;
    END
  END m0_wbd_dat_o[26]
  PIN m0_wbd_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 -4.000 68.910 4.000 ;
    END
  END m0_wbd_dat_o[27]
  PIN m0_wbd_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 -4.000 67.990 4.000 ;
    END
  END m0_wbd_dat_o[28]
  PIN m0_wbd_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 -4.000 67.070 4.000 ;
    END
  END m0_wbd_dat_o[29]
  PIN m0_wbd_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 -4.000 91.910 4.000 ;
    END
  END m0_wbd_dat_o[2]
  PIN m0_wbd_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 -4.000 66.150 4.000 ;
    END
  END m0_wbd_dat_o[30]
  PIN m0_wbd_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 -4.000 65.230 4.000 ;
    END
  END m0_wbd_dat_o[31]
  PIN m0_wbd_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 -4.000 90.990 4.000 ;
    END
  END m0_wbd_dat_o[3]
  PIN m0_wbd_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 -4.000 90.070 4.000 ;
    END
  END m0_wbd_dat_o[4]
  PIN m0_wbd_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 -4.000 89.150 4.000 ;
    END
  END m0_wbd_dat_o[5]
  PIN m0_wbd_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 -4.000 88.230 4.000 ;
    END
  END m0_wbd_dat_o[6]
  PIN m0_wbd_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 -4.000 87.310 4.000 ;
    END
  END m0_wbd_dat_o[7]
  PIN m0_wbd_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 -4.000 86.390 4.000 ;
    END
  END m0_wbd_dat_o[8]
  PIN m0_wbd_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 -4.000 85.470 4.000 ;
    END
  END m0_wbd_dat_o[9]
  PIN m0_wbd_err_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 -4.000 95.590 4.000 ;
    END
  END m0_wbd_err_o
  PIN m0_wbd_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 -4.000 34.870 4.000 ;
    END
  END m0_wbd_sel_i[0]
  PIN m0_wbd_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 -4.000 33.950 4.000 ;
    END
  END m0_wbd_sel_i[1]
  PIN m0_wbd_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 -4.000 33.030 4.000 ;
    END
  END m0_wbd_sel_i[2]
  PIN m0_wbd_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 -4.000 32.110 4.000 ;
    END
  END m0_wbd_sel_i[3]
  PIN m0_wbd_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 -4.000 0.830 4.000 ;
    END
  END m0_wbd_stb_i
  PIN m0_wbd_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 -4.000 1.750 4.000 ;
    END
  END m0_wbd_we_i
  PIN m1_wbd_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 -4.000 294.310 4.000 ;
    END
  END m1_wbd_ack_o
  PIN m1_wbd_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 -4.000 230.830 4.000 ;
    END
  END m1_wbd_adr_i[0]
  PIN m1_wbd_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 -4.000 221.630 4.000 ;
    END
  END m1_wbd_adr_i[10]
  PIN m1_wbd_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 -4.000 220.710 4.000 ;
    END
  END m1_wbd_adr_i[11]
  PIN m1_wbd_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 -4.000 219.790 4.000 ;
    END
  END m1_wbd_adr_i[12]
  PIN m1_wbd_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 -4.000 218.870 4.000 ;
    END
  END m1_wbd_adr_i[13]
  PIN m1_wbd_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 -4.000 217.950 4.000 ;
    END
  END m1_wbd_adr_i[14]
  PIN m1_wbd_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 -4.000 217.030 4.000 ;
    END
  END m1_wbd_adr_i[15]
  PIN m1_wbd_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 -4.000 216.110 4.000 ;
    END
  END m1_wbd_adr_i[16]
  PIN m1_wbd_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 -4.000 215.190 4.000 ;
    END
  END m1_wbd_adr_i[17]
  PIN m1_wbd_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 -4.000 214.270 4.000 ;
    END
  END m1_wbd_adr_i[18]
  PIN m1_wbd_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 -4.000 213.350 4.000 ;
    END
  END m1_wbd_adr_i[19]
  PIN m1_wbd_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 -4.000 229.910 4.000 ;
    END
  END m1_wbd_adr_i[1]
  PIN m1_wbd_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 -4.000 212.430 4.000 ;
    END
  END m1_wbd_adr_i[20]
  PIN m1_wbd_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 -4.000 211.510 4.000 ;
    END
  END m1_wbd_adr_i[21]
  PIN m1_wbd_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 -4.000 210.590 4.000 ;
    END
  END m1_wbd_adr_i[22]
  PIN m1_wbd_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 -4.000 209.670 4.000 ;
    END
  END m1_wbd_adr_i[23]
  PIN m1_wbd_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 -4.000 208.750 4.000 ;
    END
  END m1_wbd_adr_i[24]
  PIN m1_wbd_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 -4.000 207.830 4.000 ;
    END
  END m1_wbd_adr_i[25]
  PIN m1_wbd_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 -4.000 206.910 4.000 ;
    END
  END m1_wbd_adr_i[26]
  PIN m1_wbd_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 -4.000 205.990 4.000 ;
    END
  END m1_wbd_adr_i[27]
  PIN m1_wbd_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 -4.000 205.070 4.000 ;
    END
  END m1_wbd_adr_i[28]
  PIN m1_wbd_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 -4.000 204.150 4.000 ;
    END
  END m1_wbd_adr_i[29]
  PIN m1_wbd_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 -4.000 228.990 4.000 ;
    END
  END m1_wbd_adr_i[2]
  PIN m1_wbd_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 -4.000 203.230 4.000 ;
    END
  END m1_wbd_adr_i[30]
  PIN m1_wbd_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 -4.000 202.310 4.000 ;
    END
  END m1_wbd_adr_i[31]
  PIN m1_wbd_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 -4.000 228.070 4.000 ;
    END
  END m1_wbd_adr_i[3]
  PIN m1_wbd_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 -4.000 227.150 4.000 ;
    END
  END m1_wbd_adr_i[4]
  PIN m1_wbd_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 -4.000 226.230 4.000 ;
    END
  END m1_wbd_adr_i[5]
  PIN m1_wbd_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 -4.000 225.310 4.000 ;
    END
  END m1_wbd_adr_i[6]
  PIN m1_wbd_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 -4.000 224.390 4.000 ;
    END
  END m1_wbd_adr_i[7]
  PIN m1_wbd_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 -4.000 223.470 4.000 ;
    END
  END m1_wbd_adr_i[8]
  PIN m1_wbd_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 -4.000 222.550 4.000 ;
    END
  END m1_wbd_adr_i[9]
  PIN m1_wbd_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 -4.000 296.150 4.000 ;
    END
  END m1_wbd_cyc_i
  PIN m1_wbd_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 -4.000 263.950 4.000 ;
    END
  END m1_wbd_dat_i[0]
  PIN m1_wbd_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 -4.000 254.750 4.000 ;
    END
  END m1_wbd_dat_i[10]
  PIN m1_wbd_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 -4.000 253.830 4.000 ;
    END
  END m1_wbd_dat_i[11]
  PIN m1_wbd_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 -4.000 252.910 4.000 ;
    END
  END m1_wbd_dat_i[12]
  PIN m1_wbd_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 -4.000 251.990 4.000 ;
    END
  END m1_wbd_dat_i[13]
  PIN m1_wbd_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 -4.000 251.070 4.000 ;
    END
  END m1_wbd_dat_i[14]
  PIN m1_wbd_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 -4.000 250.150 4.000 ;
    END
  END m1_wbd_dat_i[15]
  PIN m1_wbd_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 -4.000 249.230 4.000 ;
    END
  END m1_wbd_dat_i[16]
  PIN m1_wbd_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 -4.000 248.310 4.000 ;
    END
  END m1_wbd_dat_i[17]
  PIN m1_wbd_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 -4.000 247.390 4.000 ;
    END
  END m1_wbd_dat_i[18]
  PIN m1_wbd_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 -4.000 246.470 4.000 ;
    END
  END m1_wbd_dat_i[19]
  PIN m1_wbd_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 -4.000 263.030 4.000 ;
    END
  END m1_wbd_dat_i[1]
  PIN m1_wbd_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 -4.000 245.550 4.000 ;
    END
  END m1_wbd_dat_i[20]
  PIN m1_wbd_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 -4.000 244.630 4.000 ;
    END
  END m1_wbd_dat_i[21]
  PIN m1_wbd_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 -4.000 243.710 4.000 ;
    END
  END m1_wbd_dat_i[22]
  PIN m1_wbd_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 -4.000 242.790 4.000 ;
    END
  END m1_wbd_dat_i[23]
  PIN m1_wbd_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 -4.000 241.870 4.000 ;
    END
  END m1_wbd_dat_i[24]
  PIN m1_wbd_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 -4.000 240.950 4.000 ;
    END
  END m1_wbd_dat_i[25]
  PIN m1_wbd_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 -4.000 240.030 4.000 ;
    END
  END m1_wbd_dat_i[26]
  PIN m1_wbd_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 -4.000 239.110 4.000 ;
    END
  END m1_wbd_dat_i[27]
  PIN m1_wbd_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 -4.000 238.190 4.000 ;
    END
  END m1_wbd_dat_i[28]
  PIN m1_wbd_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 -4.000 237.270 4.000 ;
    END
  END m1_wbd_dat_i[29]
  PIN m1_wbd_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 -4.000 262.110 4.000 ;
    END
  END m1_wbd_dat_i[2]
  PIN m1_wbd_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 -4.000 236.350 4.000 ;
    END
  END m1_wbd_dat_i[30]
  PIN m1_wbd_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 -4.000 235.430 4.000 ;
    END
  END m1_wbd_dat_i[31]
  PIN m1_wbd_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 -4.000 261.190 4.000 ;
    END
  END m1_wbd_dat_i[3]
  PIN m1_wbd_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 -4.000 260.270 4.000 ;
    END
  END m1_wbd_dat_i[4]
  PIN m1_wbd_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 -4.000 259.350 4.000 ;
    END
  END m1_wbd_dat_i[5]
  PIN m1_wbd_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 -4.000 258.430 4.000 ;
    END
  END m1_wbd_dat_i[6]
  PIN m1_wbd_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 -4.000 257.510 4.000 ;
    END
  END m1_wbd_dat_i[7]
  PIN m1_wbd_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 -4.000 256.590 4.000 ;
    END
  END m1_wbd_dat_i[8]
  PIN m1_wbd_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 -4.000 255.670 4.000 ;
    END
  END m1_wbd_dat_i[9]
  PIN m1_wbd_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 -4.000 293.390 4.000 ;
    END
  END m1_wbd_dat_o[0]
  PIN m1_wbd_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 -4.000 284.190 4.000 ;
    END
  END m1_wbd_dat_o[10]
  PIN m1_wbd_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 -4.000 283.270 4.000 ;
    END
  END m1_wbd_dat_o[11]
  PIN m1_wbd_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 -4.000 282.350 4.000 ;
    END
  END m1_wbd_dat_o[12]
  PIN m1_wbd_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 -4.000 281.430 4.000 ;
    END
  END m1_wbd_dat_o[13]
  PIN m1_wbd_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 -4.000 280.510 4.000 ;
    END
  END m1_wbd_dat_o[14]
  PIN m1_wbd_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 -4.000 279.590 4.000 ;
    END
  END m1_wbd_dat_o[15]
  PIN m1_wbd_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 -4.000 278.670 4.000 ;
    END
  END m1_wbd_dat_o[16]
  PIN m1_wbd_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 -4.000 277.750 4.000 ;
    END
  END m1_wbd_dat_o[17]
  PIN m1_wbd_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 -4.000 276.830 4.000 ;
    END
  END m1_wbd_dat_o[18]
  PIN m1_wbd_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 -4.000 275.910 4.000 ;
    END
  END m1_wbd_dat_o[19]
  PIN m1_wbd_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 -4.000 292.470 4.000 ;
    END
  END m1_wbd_dat_o[1]
  PIN m1_wbd_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 -4.000 274.990 4.000 ;
    END
  END m1_wbd_dat_o[20]
  PIN m1_wbd_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 -4.000 274.070 4.000 ;
    END
  END m1_wbd_dat_o[21]
  PIN m1_wbd_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 -4.000 273.150 4.000 ;
    END
  END m1_wbd_dat_o[22]
  PIN m1_wbd_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 -4.000 272.230 4.000 ;
    END
  END m1_wbd_dat_o[23]
  PIN m1_wbd_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 -4.000 271.310 4.000 ;
    END
  END m1_wbd_dat_o[24]
  PIN m1_wbd_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 -4.000 270.390 4.000 ;
    END
  END m1_wbd_dat_o[25]
  PIN m1_wbd_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 -4.000 269.470 4.000 ;
    END
  END m1_wbd_dat_o[26]
  PIN m1_wbd_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 -4.000 268.550 4.000 ;
    END
  END m1_wbd_dat_o[27]
  PIN m1_wbd_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 -4.000 267.630 4.000 ;
    END
  END m1_wbd_dat_o[28]
  PIN m1_wbd_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 -4.000 266.710 4.000 ;
    END
  END m1_wbd_dat_o[29]
  PIN m1_wbd_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 -4.000 291.550 4.000 ;
    END
  END m1_wbd_dat_o[2]
  PIN m1_wbd_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 -4.000 265.790 4.000 ;
    END
  END m1_wbd_dat_o[30]
  PIN m1_wbd_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 -4.000 264.870 4.000 ;
    END
  END m1_wbd_dat_o[31]
  PIN m1_wbd_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 -4.000 290.630 4.000 ;
    END
  END m1_wbd_dat_o[3]
  PIN m1_wbd_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 -4.000 289.710 4.000 ;
    END
  END m1_wbd_dat_o[4]
  PIN m1_wbd_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 -4.000 288.790 4.000 ;
    END
  END m1_wbd_dat_o[5]
  PIN m1_wbd_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 -4.000 287.870 4.000 ;
    END
  END m1_wbd_dat_o[6]
  PIN m1_wbd_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 -4.000 286.950 4.000 ;
    END
  END m1_wbd_dat_o[7]
  PIN m1_wbd_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 -4.000 286.030 4.000 ;
    END
  END m1_wbd_dat_o[8]
  PIN m1_wbd_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 -4.000 285.110 4.000 ;
    END
  END m1_wbd_dat_o[9]
  PIN m1_wbd_err_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 -4.000 295.230 4.000 ;
    END
  END m1_wbd_err_o
  PIN m1_wbd_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 -4.000 234.510 4.000 ;
    END
  END m1_wbd_sel_i[0]
  PIN m1_wbd_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 -4.000 233.590 4.000 ;
    END
  END m1_wbd_sel_i[1]
  PIN m1_wbd_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 -4.000 232.670 4.000 ;
    END
  END m1_wbd_sel_i[2]
  PIN m1_wbd_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 -4.000 231.750 4.000 ;
    END
  END m1_wbd_sel_i[3]
  PIN m1_wbd_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 -4.000 200.470 4.000 ;
    END
  END m1_wbd_stb_i
  PIN m1_wbd_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 -4.000 201.390 4.000 ;
    END
  END m1_wbd_we_i
  PIN m2_wbd_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 -4.000 794.330 4.000 ;
    END
  END m2_wbd_ack_o
  PIN m2_wbd_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 -4.000 730.850 4.000 ;
    END
  END m2_wbd_adr_i[0]
  PIN m2_wbd_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 -4.000 721.650 4.000 ;
    END
  END m2_wbd_adr_i[10]
  PIN m2_wbd_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 -4.000 720.730 4.000 ;
    END
  END m2_wbd_adr_i[11]
  PIN m2_wbd_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 -4.000 719.810 4.000 ;
    END
  END m2_wbd_adr_i[12]
  PIN m2_wbd_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 -4.000 718.890 4.000 ;
    END
  END m2_wbd_adr_i[13]
  PIN m2_wbd_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 -4.000 717.970 4.000 ;
    END
  END m2_wbd_adr_i[14]
  PIN m2_wbd_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 -4.000 717.050 4.000 ;
    END
  END m2_wbd_adr_i[15]
  PIN m2_wbd_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 -4.000 716.130 4.000 ;
    END
  END m2_wbd_adr_i[16]
  PIN m2_wbd_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 -4.000 715.210 4.000 ;
    END
  END m2_wbd_adr_i[17]
  PIN m2_wbd_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 -4.000 714.290 4.000 ;
    END
  END m2_wbd_adr_i[18]
  PIN m2_wbd_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 -4.000 713.370 4.000 ;
    END
  END m2_wbd_adr_i[19]
  PIN m2_wbd_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 -4.000 729.930 4.000 ;
    END
  END m2_wbd_adr_i[1]
  PIN m2_wbd_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 -4.000 712.450 4.000 ;
    END
  END m2_wbd_adr_i[20]
  PIN m2_wbd_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 -4.000 711.530 4.000 ;
    END
  END m2_wbd_adr_i[21]
  PIN m2_wbd_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 -4.000 710.610 4.000 ;
    END
  END m2_wbd_adr_i[22]
  PIN m2_wbd_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 -4.000 709.690 4.000 ;
    END
  END m2_wbd_adr_i[23]
  PIN m2_wbd_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 -4.000 708.770 4.000 ;
    END
  END m2_wbd_adr_i[24]
  PIN m2_wbd_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 -4.000 707.850 4.000 ;
    END
  END m2_wbd_adr_i[25]
  PIN m2_wbd_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 -4.000 706.930 4.000 ;
    END
  END m2_wbd_adr_i[26]
  PIN m2_wbd_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 -4.000 706.010 4.000 ;
    END
  END m2_wbd_adr_i[27]
  PIN m2_wbd_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 -4.000 705.090 4.000 ;
    END
  END m2_wbd_adr_i[28]
  PIN m2_wbd_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 -4.000 704.170 4.000 ;
    END
  END m2_wbd_adr_i[29]
  PIN m2_wbd_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 -4.000 729.010 4.000 ;
    END
  END m2_wbd_adr_i[2]
  PIN m2_wbd_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.970 -4.000 703.250 4.000 ;
    END
  END m2_wbd_adr_i[30]
  PIN m2_wbd_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 -4.000 702.330 4.000 ;
    END
  END m2_wbd_adr_i[31]
  PIN m2_wbd_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 -4.000 728.090 4.000 ;
    END
  END m2_wbd_adr_i[3]
  PIN m2_wbd_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 -4.000 727.170 4.000 ;
    END
  END m2_wbd_adr_i[4]
  PIN m2_wbd_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.970 -4.000 726.250 4.000 ;
    END
  END m2_wbd_adr_i[5]
  PIN m2_wbd_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 -4.000 725.330 4.000 ;
    END
  END m2_wbd_adr_i[6]
  PIN m2_wbd_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 -4.000 724.410 4.000 ;
    END
  END m2_wbd_adr_i[7]
  PIN m2_wbd_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 -4.000 723.490 4.000 ;
    END
  END m2_wbd_adr_i[8]
  PIN m2_wbd_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 -4.000 722.570 4.000 ;
    END
  END m2_wbd_adr_i[9]
  PIN m2_wbd_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 -4.000 796.170 4.000 ;
    END
  END m2_wbd_cyc_i
  PIN m2_wbd_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 -4.000 763.970 4.000 ;
    END
  END m2_wbd_dat_i[0]
  PIN m2_wbd_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 -4.000 754.770 4.000 ;
    END
  END m2_wbd_dat_i[10]
  PIN m2_wbd_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 -4.000 753.850 4.000 ;
    END
  END m2_wbd_dat_i[11]
  PIN m2_wbd_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 -4.000 752.930 4.000 ;
    END
  END m2_wbd_dat_i[12]
  PIN m2_wbd_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.730 -4.000 752.010 4.000 ;
    END
  END m2_wbd_dat_i[13]
  PIN m2_wbd_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 -4.000 751.090 4.000 ;
    END
  END m2_wbd_dat_i[14]
  PIN m2_wbd_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 -4.000 750.170 4.000 ;
    END
  END m2_wbd_dat_i[15]
  PIN m2_wbd_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 -4.000 749.250 4.000 ;
    END
  END m2_wbd_dat_i[16]
  PIN m2_wbd_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 -4.000 748.330 4.000 ;
    END
  END m2_wbd_dat_i[17]
  PIN m2_wbd_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 -4.000 747.410 4.000 ;
    END
  END m2_wbd_dat_i[18]
  PIN m2_wbd_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 -4.000 746.490 4.000 ;
    END
  END m2_wbd_dat_i[19]
  PIN m2_wbd_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.770 -4.000 763.050 4.000 ;
    END
  END m2_wbd_dat_i[1]
  PIN m2_wbd_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 -4.000 745.570 4.000 ;
    END
  END m2_wbd_dat_i[20]
  PIN m2_wbd_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.370 -4.000 744.650 4.000 ;
    END
  END m2_wbd_dat_i[21]
  PIN m2_wbd_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 -4.000 743.730 4.000 ;
    END
  END m2_wbd_dat_i[22]
  PIN m2_wbd_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 -4.000 742.810 4.000 ;
    END
  END m2_wbd_dat_i[23]
  PIN m2_wbd_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 -4.000 741.890 4.000 ;
    END
  END m2_wbd_dat_i[24]
  PIN m2_wbd_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 -4.000 740.970 4.000 ;
    END
  END m2_wbd_dat_i[25]
  PIN m2_wbd_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 -4.000 740.050 4.000 ;
    END
  END m2_wbd_dat_i[26]
  PIN m2_wbd_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.850 -4.000 739.130 4.000 ;
    END
  END m2_wbd_dat_i[27]
  PIN m2_wbd_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 -4.000 738.210 4.000 ;
    END
  END m2_wbd_dat_i[28]
  PIN m2_wbd_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 -4.000 737.290 4.000 ;
    END
  END m2_wbd_dat_i[29]
  PIN m2_wbd_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.850 -4.000 762.130 4.000 ;
    END
  END m2_wbd_dat_i[2]
  PIN m2_wbd_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.090 -4.000 736.370 4.000 ;
    END
  END m2_wbd_dat_i[30]
  PIN m2_wbd_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 -4.000 735.450 4.000 ;
    END
  END m2_wbd_dat_i[31]
  PIN m2_wbd_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930 -4.000 761.210 4.000 ;
    END
  END m2_wbd_dat_i[3]
  PIN m2_wbd_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 -4.000 760.290 4.000 ;
    END
  END m2_wbd_dat_i[4]
  PIN m2_wbd_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 -4.000 759.370 4.000 ;
    END
  END m2_wbd_dat_i[5]
  PIN m2_wbd_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 -4.000 758.450 4.000 ;
    END
  END m2_wbd_dat_i[6]
  PIN m2_wbd_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 -4.000 757.530 4.000 ;
    END
  END m2_wbd_dat_i[7]
  PIN m2_wbd_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.330 -4.000 756.610 4.000 ;
    END
  END m2_wbd_dat_i[8]
  PIN m2_wbd_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.410 -4.000 755.690 4.000 ;
    END
  END m2_wbd_dat_i[9]
  PIN m2_wbd_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 -4.000 793.410 4.000 ;
    END
  END m2_wbd_dat_o[0]
  PIN m2_wbd_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 -4.000 784.210 4.000 ;
    END
  END m2_wbd_dat_o[10]
  PIN m2_wbd_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 -4.000 783.290 4.000 ;
    END
  END m2_wbd_dat_o[11]
  PIN m2_wbd_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 -4.000 782.370 4.000 ;
    END
  END m2_wbd_dat_o[12]
  PIN m2_wbd_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 -4.000 781.450 4.000 ;
    END
  END m2_wbd_dat_o[13]
  PIN m2_wbd_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 -4.000 780.530 4.000 ;
    END
  END m2_wbd_dat_o[14]
  PIN m2_wbd_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 -4.000 779.610 4.000 ;
    END
  END m2_wbd_dat_o[15]
  PIN m2_wbd_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 -4.000 778.690 4.000 ;
    END
  END m2_wbd_dat_o[16]
  PIN m2_wbd_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 -4.000 777.770 4.000 ;
    END
  END m2_wbd_dat_o[17]
  PIN m2_wbd_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 -4.000 776.850 4.000 ;
    END
  END m2_wbd_dat_o[18]
  PIN m2_wbd_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 -4.000 775.930 4.000 ;
    END
  END m2_wbd_dat_o[19]
  PIN m2_wbd_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 -4.000 792.490 4.000 ;
    END
  END m2_wbd_dat_o[1]
  PIN m2_wbd_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 -4.000 775.010 4.000 ;
    END
  END m2_wbd_dat_o[20]
  PIN m2_wbd_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.810 -4.000 774.090 4.000 ;
    END
  END m2_wbd_dat_o[21]
  PIN m2_wbd_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 -4.000 773.170 4.000 ;
    END
  END m2_wbd_dat_o[22]
  PIN m2_wbd_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 -4.000 772.250 4.000 ;
    END
  END m2_wbd_dat_o[23]
  PIN m2_wbd_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.050 -4.000 771.330 4.000 ;
    END
  END m2_wbd_dat_o[24]
  PIN m2_wbd_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 -4.000 770.410 4.000 ;
    END
  END m2_wbd_dat_o[25]
  PIN m2_wbd_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.210 -4.000 769.490 4.000 ;
    END
  END m2_wbd_dat_o[26]
  PIN m2_wbd_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.290 -4.000 768.570 4.000 ;
    END
  END m2_wbd_dat_o[27]
  PIN m2_wbd_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 -4.000 767.650 4.000 ;
    END
  END m2_wbd_dat_o[28]
  PIN m2_wbd_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 -4.000 766.730 4.000 ;
    END
  END m2_wbd_dat_o[29]
  PIN m2_wbd_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 -4.000 791.570 4.000 ;
    END
  END m2_wbd_dat_o[2]
  PIN m2_wbd_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 -4.000 765.810 4.000 ;
    END
  END m2_wbd_dat_o[30]
  PIN m2_wbd_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 -4.000 764.890 4.000 ;
    END
  END m2_wbd_dat_o[31]
  PIN m2_wbd_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.370 -4.000 790.650 4.000 ;
    END
  END m2_wbd_dat_o[3]
  PIN m2_wbd_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 -4.000 789.730 4.000 ;
    END
  END m2_wbd_dat_o[4]
  PIN m2_wbd_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.530 -4.000 788.810 4.000 ;
    END
  END m2_wbd_dat_o[5]
  PIN m2_wbd_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.610 -4.000 787.890 4.000 ;
    END
  END m2_wbd_dat_o[6]
  PIN m2_wbd_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 -4.000 786.970 4.000 ;
    END
  END m2_wbd_dat_o[7]
  PIN m2_wbd_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 -4.000 786.050 4.000 ;
    END
  END m2_wbd_dat_o[8]
  PIN m2_wbd_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 -4.000 785.130 4.000 ;
    END
  END m2_wbd_dat_o[9]
  PIN m2_wbd_err_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.970 -4.000 795.250 4.000 ;
    END
  END m2_wbd_err_o
  PIN m2_wbd_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 -4.000 734.530 4.000 ;
    END
  END m2_wbd_sel_i[0]
  PIN m2_wbd_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 -4.000 733.610 4.000 ;
    END
  END m2_wbd_sel_i[1]
  PIN m2_wbd_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 -4.000 732.690 4.000 ;
    END
  END m2_wbd_sel_i[2]
  PIN m2_wbd_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 -4.000 731.770 4.000 ;
    END
  END m2_wbd_sel_i[3]
  PIN m2_wbd_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 -4.000 700.490 4.000 ;
    END
  END m2_wbd_stb_i
  PIN m2_wbd_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 -4.000 701.410 4.000 ;
    END
  END m2_wbd_we_i
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2196.000 2.080 2204.000 2.680 ;
    END
  END rst_n
  PIN s0_wbd_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 146.000 94.670 154.000 ;
    END
  END s0_wbd_ack_i
  PIN s0_wbd_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 146.000 31.190 154.000 ;
    END
  END s0_wbd_adr_o[0]
  PIN s0_wbd_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 146.000 21.990 154.000 ;
    END
  END s0_wbd_adr_o[10]
  PIN s0_wbd_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 146.000 21.070 154.000 ;
    END
  END s0_wbd_adr_o[11]
  PIN s0_wbd_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 146.000 20.150 154.000 ;
    END
  END s0_wbd_adr_o[12]
  PIN s0_wbd_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 146.000 19.230 154.000 ;
    END
  END s0_wbd_adr_o[13]
  PIN s0_wbd_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 146.000 18.310 154.000 ;
    END
  END s0_wbd_adr_o[14]
  PIN s0_wbd_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 146.000 17.390 154.000 ;
    END
  END s0_wbd_adr_o[15]
  PIN s0_wbd_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 146.000 16.470 154.000 ;
    END
  END s0_wbd_adr_o[16]
  PIN s0_wbd_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 146.000 15.550 154.000 ;
    END
  END s0_wbd_adr_o[17]
  PIN s0_wbd_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 146.000 14.630 154.000 ;
    END
  END s0_wbd_adr_o[18]
  PIN s0_wbd_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 146.000 13.710 154.000 ;
    END
  END s0_wbd_adr_o[19]
  PIN s0_wbd_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 146.000 30.270 154.000 ;
    END
  END s0_wbd_adr_o[1]
  PIN s0_wbd_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 146.000 12.790 154.000 ;
    END
  END s0_wbd_adr_o[20]
  PIN s0_wbd_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 146.000 11.870 154.000 ;
    END
  END s0_wbd_adr_o[21]
  PIN s0_wbd_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 146.000 10.950 154.000 ;
    END
  END s0_wbd_adr_o[22]
  PIN s0_wbd_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 146.000 10.030 154.000 ;
    END
  END s0_wbd_adr_o[23]
  PIN s0_wbd_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 146.000 9.110 154.000 ;
    END
  END s0_wbd_adr_o[24]
  PIN s0_wbd_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 146.000 8.190 154.000 ;
    END
  END s0_wbd_adr_o[25]
  PIN s0_wbd_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 146.000 7.270 154.000 ;
    END
  END s0_wbd_adr_o[26]
  PIN s0_wbd_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 146.000 6.350 154.000 ;
    END
  END s0_wbd_adr_o[27]
  PIN s0_wbd_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 146.000 5.430 154.000 ;
    END
  END s0_wbd_adr_o[28]
  PIN s0_wbd_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 146.000 4.510 154.000 ;
    END
  END s0_wbd_adr_o[29]
  PIN s0_wbd_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 146.000 29.350 154.000 ;
    END
  END s0_wbd_adr_o[2]
  PIN s0_wbd_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 146.000 3.590 154.000 ;
    END
  END s0_wbd_adr_o[30]
  PIN s0_wbd_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 146.000 2.670 154.000 ;
    END
  END s0_wbd_adr_o[31]
  PIN s0_wbd_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 146.000 28.430 154.000 ;
    END
  END s0_wbd_adr_o[3]
  PIN s0_wbd_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 146.000 27.510 154.000 ;
    END
  END s0_wbd_adr_o[4]
  PIN s0_wbd_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 146.000 26.590 154.000 ;
    END
  END s0_wbd_adr_o[5]
  PIN s0_wbd_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 146.000 25.670 154.000 ;
    END
  END s0_wbd_adr_o[6]
  PIN s0_wbd_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 146.000 24.750 154.000 ;
    END
  END s0_wbd_adr_o[7]
  PIN s0_wbd_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 146.000 23.830 154.000 ;
    END
  END s0_wbd_adr_o[8]
  PIN s0_wbd_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 146.000 22.910 154.000 ;
    END
  END s0_wbd_adr_o[9]
  PIN s0_wbd_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 146.000 95.590 154.000 ;
    END
  END s0_wbd_cyc_o
  PIN s0_wbd_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 146.000 93.750 154.000 ;
    END
  END s0_wbd_dat_i[0]
  PIN s0_wbd_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 146.000 84.550 154.000 ;
    END
  END s0_wbd_dat_i[10]
  PIN s0_wbd_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 146.000 83.630 154.000 ;
    END
  END s0_wbd_dat_i[11]
  PIN s0_wbd_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 146.000 82.710 154.000 ;
    END
  END s0_wbd_dat_i[12]
  PIN s0_wbd_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 146.000 81.790 154.000 ;
    END
  END s0_wbd_dat_i[13]
  PIN s0_wbd_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 146.000 80.870 154.000 ;
    END
  END s0_wbd_dat_i[14]
  PIN s0_wbd_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 146.000 79.950 154.000 ;
    END
  END s0_wbd_dat_i[15]
  PIN s0_wbd_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 146.000 79.030 154.000 ;
    END
  END s0_wbd_dat_i[16]
  PIN s0_wbd_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 146.000 78.110 154.000 ;
    END
  END s0_wbd_dat_i[17]
  PIN s0_wbd_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 146.000 77.190 154.000 ;
    END
  END s0_wbd_dat_i[18]
  PIN s0_wbd_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 146.000 76.270 154.000 ;
    END
  END s0_wbd_dat_i[19]
  PIN s0_wbd_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 146.000 92.830 154.000 ;
    END
  END s0_wbd_dat_i[1]
  PIN s0_wbd_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 146.000 75.350 154.000 ;
    END
  END s0_wbd_dat_i[20]
  PIN s0_wbd_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 146.000 74.430 154.000 ;
    END
  END s0_wbd_dat_i[21]
  PIN s0_wbd_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 146.000 73.510 154.000 ;
    END
  END s0_wbd_dat_i[22]
  PIN s0_wbd_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 146.000 72.590 154.000 ;
    END
  END s0_wbd_dat_i[23]
  PIN s0_wbd_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 146.000 71.670 154.000 ;
    END
  END s0_wbd_dat_i[24]
  PIN s0_wbd_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 146.000 70.750 154.000 ;
    END
  END s0_wbd_dat_i[25]
  PIN s0_wbd_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 146.000 69.830 154.000 ;
    END
  END s0_wbd_dat_i[26]
  PIN s0_wbd_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 146.000 68.910 154.000 ;
    END
  END s0_wbd_dat_i[27]
  PIN s0_wbd_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 146.000 67.990 154.000 ;
    END
  END s0_wbd_dat_i[28]
  PIN s0_wbd_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 146.000 67.070 154.000 ;
    END
  END s0_wbd_dat_i[29]
  PIN s0_wbd_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 146.000 91.910 154.000 ;
    END
  END s0_wbd_dat_i[2]
  PIN s0_wbd_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 146.000 66.150 154.000 ;
    END
  END s0_wbd_dat_i[30]
  PIN s0_wbd_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 146.000 65.230 154.000 ;
    END
  END s0_wbd_dat_i[31]
  PIN s0_wbd_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 146.000 90.990 154.000 ;
    END
  END s0_wbd_dat_i[3]
  PIN s0_wbd_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 146.000 90.070 154.000 ;
    END
  END s0_wbd_dat_i[4]
  PIN s0_wbd_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 146.000 89.150 154.000 ;
    END
  END s0_wbd_dat_i[5]
  PIN s0_wbd_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 146.000 88.230 154.000 ;
    END
  END s0_wbd_dat_i[6]
  PIN s0_wbd_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 146.000 87.310 154.000 ;
    END
  END s0_wbd_dat_i[7]
  PIN s0_wbd_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 146.000 86.390 154.000 ;
    END
  END s0_wbd_dat_i[8]
  PIN s0_wbd_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 146.000 85.470 154.000 ;
    END
  END s0_wbd_dat_i[9]
  PIN s0_wbd_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 146.000 64.310 154.000 ;
    END
  END s0_wbd_dat_o[0]
  PIN s0_wbd_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 146.000 55.110 154.000 ;
    END
  END s0_wbd_dat_o[10]
  PIN s0_wbd_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 146.000 54.190 154.000 ;
    END
  END s0_wbd_dat_o[11]
  PIN s0_wbd_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 146.000 53.270 154.000 ;
    END
  END s0_wbd_dat_o[12]
  PIN s0_wbd_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 146.000 52.350 154.000 ;
    END
  END s0_wbd_dat_o[13]
  PIN s0_wbd_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 146.000 51.430 154.000 ;
    END
  END s0_wbd_dat_o[14]
  PIN s0_wbd_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 146.000 50.510 154.000 ;
    END
  END s0_wbd_dat_o[15]
  PIN s0_wbd_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 146.000 49.590 154.000 ;
    END
  END s0_wbd_dat_o[16]
  PIN s0_wbd_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 146.000 48.670 154.000 ;
    END
  END s0_wbd_dat_o[17]
  PIN s0_wbd_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 146.000 47.750 154.000 ;
    END
  END s0_wbd_dat_o[18]
  PIN s0_wbd_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 146.000 46.830 154.000 ;
    END
  END s0_wbd_dat_o[19]
  PIN s0_wbd_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 146.000 63.390 154.000 ;
    END
  END s0_wbd_dat_o[1]
  PIN s0_wbd_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 146.000 45.910 154.000 ;
    END
  END s0_wbd_dat_o[20]
  PIN s0_wbd_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 146.000 44.990 154.000 ;
    END
  END s0_wbd_dat_o[21]
  PIN s0_wbd_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 146.000 44.070 154.000 ;
    END
  END s0_wbd_dat_o[22]
  PIN s0_wbd_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 146.000 43.150 154.000 ;
    END
  END s0_wbd_dat_o[23]
  PIN s0_wbd_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 146.000 42.230 154.000 ;
    END
  END s0_wbd_dat_o[24]
  PIN s0_wbd_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 146.000 41.310 154.000 ;
    END
  END s0_wbd_dat_o[25]
  PIN s0_wbd_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 146.000 40.390 154.000 ;
    END
  END s0_wbd_dat_o[26]
  PIN s0_wbd_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 146.000 39.470 154.000 ;
    END
  END s0_wbd_dat_o[27]
  PIN s0_wbd_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 146.000 38.550 154.000 ;
    END
  END s0_wbd_dat_o[28]
  PIN s0_wbd_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 146.000 37.630 154.000 ;
    END
  END s0_wbd_dat_o[29]
  PIN s0_wbd_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 146.000 62.470 154.000 ;
    END
  END s0_wbd_dat_o[2]
  PIN s0_wbd_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 146.000 36.710 154.000 ;
    END
  END s0_wbd_dat_o[30]
  PIN s0_wbd_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 146.000 35.790 154.000 ;
    END
  END s0_wbd_dat_o[31]
  PIN s0_wbd_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 146.000 61.550 154.000 ;
    END
  END s0_wbd_dat_o[3]
  PIN s0_wbd_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 146.000 60.630 154.000 ;
    END
  END s0_wbd_dat_o[4]
  PIN s0_wbd_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 146.000 59.710 154.000 ;
    END
  END s0_wbd_dat_o[5]
  PIN s0_wbd_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 146.000 58.790 154.000 ;
    END
  END s0_wbd_dat_o[6]
  PIN s0_wbd_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 146.000 57.870 154.000 ;
    END
  END s0_wbd_dat_o[7]
  PIN s0_wbd_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 146.000 56.950 154.000 ;
    END
  END s0_wbd_dat_o[8]
  PIN s0_wbd_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 146.000 56.030 154.000 ;
    END
  END s0_wbd_dat_o[9]
  PIN s0_wbd_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 146.000 34.870 154.000 ;
    END
  END s0_wbd_sel_o[0]
  PIN s0_wbd_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 146.000 33.950 154.000 ;
    END
  END s0_wbd_sel_o[1]
  PIN s0_wbd_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 146.000 33.030 154.000 ;
    END
  END s0_wbd_sel_o[2]
  PIN s0_wbd_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 146.000 32.110 154.000 ;
    END
  END s0_wbd_sel_o[3]
  PIN s0_wbd_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 146.000 0.830 154.000 ;
    END
  END s0_wbd_stb_o
  PIN s0_wbd_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 146.000 1.750 154.000 ;
    END
  END s0_wbd_we_o
  PIN s1_wbd_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 146.000 794.330 154.000 ;
    END
  END s1_wbd_ack_i
  PIN s1_wbd_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 146.000 730.850 154.000 ;
    END
  END s1_wbd_adr_o[0]
  PIN s1_wbd_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 146.000 721.650 154.000 ;
    END
  END s1_wbd_adr_o[10]
  PIN s1_wbd_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 146.000 720.730 154.000 ;
    END
  END s1_wbd_adr_o[11]
  PIN s1_wbd_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 146.000 719.810 154.000 ;
    END
  END s1_wbd_adr_o[12]
  PIN s1_wbd_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 146.000 718.890 154.000 ;
    END
  END s1_wbd_adr_o[13]
  PIN s1_wbd_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 146.000 717.970 154.000 ;
    END
  END s1_wbd_adr_o[14]
  PIN s1_wbd_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 146.000 717.050 154.000 ;
    END
  END s1_wbd_adr_o[15]
  PIN s1_wbd_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 146.000 716.130 154.000 ;
    END
  END s1_wbd_adr_o[16]
  PIN s1_wbd_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 146.000 715.210 154.000 ;
    END
  END s1_wbd_adr_o[17]
  PIN s1_wbd_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 146.000 714.290 154.000 ;
    END
  END s1_wbd_adr_o[18]
  PIN s1_wbd_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 146.000 713.370 154.000 ;
    END
  END s1_wbd_adr_o[19]
  PIN s1_wbd_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 146.000 729.930 154.000 ;
    END
  END s1_wbd_adr_o[1]
  PIN s1_wbd_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 146.000 712.450 154.000 ;
    END
  END s1_wbd_adr_o[20]
  PIN s1_wbd_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 146.000 711.530 154.000 ;
    END
  END s1_wbd_adr_o[21]
  PIN s1_wbd_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 146.000 710.610 154.000 ;
    END
  END s1_wbd_adr_o[22]
  PIN s1_wbd_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 146.000 709.690 154.000 ;
    END
  END s1_wbd_adr_o[23]
  PIN s1_wbd_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 146.000 708.770 154.000 ;
    END
  END s1_wbd_adr_o[24]
  PIN s1_wbd_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 146.000 707.850 154.000 ;
    END
  END s1_wbd_adr_o[25]
  PIN s1_wbd_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 146.000 706.930 154.000 ;
    END
  END s1_wbd_adr_o[26]
  PIN s1_wbd_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 146.000 706.010 154.000 ;
    END
  END s1_wbd_adr_o[27]
  PIN s1_wbd_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 146.000 705.090 154.000 ;
    END
  END s1_wbd_adr_o[28]
  PIN s1_wbd_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 146.000 704.170 154.000 ;
    END
  END s1_wbd_adr_o[29]
  PIN s1_wbd_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 146.000 729.010 154.000 ;
    END
  END s1_wbd_adr_o[2]
  PIN s1_wbd_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.970 146.000 703.250 154.000 ;
    END
  END s1_wbd_adr_o[30]
  PIN s1_wbd_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 146.000 702.330 154.000 ;
    END
  END s1_wbd_adr_o[31]
  PIN s1_wbd_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 146.000 728.090 154.000 ;
    END
  END s1_wbd_adr_o[3]
  PIN s1_wbd_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 146.000 727.170 154.000 ;
    END
  END s1_wbd_adr_o[4]
  PIN s1_wbd_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.970 146.000 726.250 154.000 ;
    END
  END s1_wbd_adr_o[5]
  PIN s1_wbd_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 146.000 725.330 154.000 ;
    END
  END s1_wbd_adr_o[6]
  PIN s1_wbd_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 146.000 724.410 154.000 ;
    END
  END s1_wbd_adr_o[7]
  PIN s1_wbd_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 146.000 723.490 154.000 ;
    END
  END s1_wbd_adr_o[8]
  PIN s1_wbd_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 146.000 722.570 154.000 ;
    END
  END s1_wbd_adr_o[9]
  PIN s1_wbd_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.970 146.000 795.250 154.000 ;
    END
  END s1_wbd_cyc_o
  PIN s1_wbd_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 146.000 793.410 154.000 ;
    END
  END s1_wbd_dat_i[0]
  PIN s1_wbd_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 146.000 784.210 154.000 ;
    END
  END s1_wbd_dat_i[10]
  PIN s1_wbd_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 146.000 783.290 154.000 ;
    END
  END s1_wbd_dat_i[11]
  PIN s1_wbd_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 146.000 782.370 154.000 ;
    END
  END s1_wbd_dat_i[12]
  PIN s1_wbd_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 146.000 781.450 154.000 ;
    END
  END s1_wbd_dat_i[13]
  PIN s1_wbd_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 146.000 780.530 154.000 ;
    END
  END s1_wbd_dat_i[14]
  PIN s1_wbd_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 146.000 779.610 154.000 ;
    END
  END s1_wbd_dat_i[15]
  PIN s1_wbd_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 146.000 778.690 154.000 ;
    END
  END s1_wbd_dat_i[16]
  PIN s1_wbd_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 146.000 777.770 154.000 ;
    END
  END s1_wbd_dat_i[17]
  PIN s1_wbd_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 146.000 776.850 154.000 ;
    END
  END s1_wbd_dat_i[18]
  PIN s1_wbd_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 146.000 775.930 154.000 ;
    END
  END s1_wbd_dat_i[19]
  PIN s1_wbd_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 146.000 792.490 154.000 ;
    END
  END s1_wbd_dat_i[1]
  PIN s1_wbd_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 146.000 775.010 154.000 ;
    END
  END s1_wbd_dat_i[20]
  PIN s1_wbd_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.810 146.000 774.090 154.000 ;
    END
  END s1_wbd_dat_i[21]
  PIN s1_wbd_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 146.000 773.170 154.000 ;
    END
  END s1_wbd_dat_i[22]
  PIN s1_wbd_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 146.000 772.250 154.000 ;
    END
  END s1_wbd_dat_i[23]
  PIN s1_wbd_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.050 146.000 771.330 154.000 ;
    END
  END s1_wbd_dat_i[24]
  PIN s1_wbd_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 146.000 770.410 154.000 ;
    END
  END s1_wbd_dat_i[25]
  PIN s1_wbd_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.210 146.000 769.490 154.000 ;
    END
  END s1_wbd_dat_i[26]
  PIN s1_wbd_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.290 146.000 768.570 154.000 ;
    END
  END s1_wbd_dat_i[27]
  PIN s1_wbd_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 146.000 767.650 154.000 ;
    END
  END s1_wbd_dat_i[28]
  PIN s1_wbd_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 146.000 766.730 154.000 ;
    END
  END s1_wbd_dat_i[29]
  PIN s1_wbd_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 146.000 791.570 154.000 ;
    END
  END s1_wbd_dat_i[2]
  PIN s1_wbd_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 146.000 765.810 154.000 ;
    END
  END s1_wbd_dat_i[30]
  PIN s1_wbd_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 146.000 764.890 154.000 ;
    END
  END s1_wbd_dat_i[31]
  PIN s1_wbd_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.370 146.000 790.650 154.000 ;
    END
  END s1_wbd_dat_i[3]
  PIN s1_wbd_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 146.000 789.730 154.000 ;
    END
  END s1_wbd_dat_i[4]
  PIN s1_wbd_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.530 146.000 788.810 154.000 ;
    END
  END s1_wbd_dat_i[5]
  PIN s1_wbd_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.610 146.000 787.890 154.000 ;
    END
  END s1_wbd_dat_i[6]
  PIN s1_wbd_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 146.000 786.970 154.000 ;
    END
  END s1_wbd_dat_i[7]
  PIN s1_wbd_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 146.000 786.050 154.000 ;
    END
  END s1_wbd_dat_i[8]
  PIN s1_wbd_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 146.000 785.130 154.000 ;
    END
  END s1_wbd_dat_i[9]
  PIN s1_wbd_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 146.000 763.970 154.000 ;
    END
  END s1_wbd_dat_o[0]
  PIN s1_wbd_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 146.000 754.770 154.000 ;
    END
  END s1_wbd_dat_o[10]
  PIN s1_wbd_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 146.000 753.850 154.000 ;
    END
  END s1_wbd_dat_o[11]
  PIN s1_wbd_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 146.000 752.930 154.000 ;
    END
  END s1_wbd_dat_o[12]
  PIN s1_wbd_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.730 146.000 752.010 154.000 ;
    END
  END s1_wbd_dat_o[13]
  PIN s1_wbd_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 146.000 751.090 154.000 ;
    END
  END s1_wbd_dat_o[14]
  PIN s1_wbd_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 146.000 750.170 154.000 ;
    END
  END s1_wbd_dat_o[15]
  PIN s1_wbd_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 146.000 749.250 154.000 ;
    END
  END s1_wbd_dat_o[16]
  PIN s1_wbd_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 146.000 748.330 154.000 ;
    END
  END s1_wbd_dat_o[17]
  PIN s1_wbd_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 146.000 747.410 154.000 ;
    END
  END s1_wbd_dat_o[18]
  PIN s1_wbd_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 146.000 746.490 154.000 ;
    END
  END s1_wbd_dat_o[19]
  PIN s1_wbd_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.770 146.000 763.050 154.000 ;
    END
  END s1_wbd_dat_o[1]
  PIN s1_wbd_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 146.000 745.570 154.000 ;
    END
  END s1_wbd_dat_o[20]
  PIN s1_wbd_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.370 146.000 744.650 154.000 ;
    END
  END s1_wbd_dat_o[21]
  PIN s1_wbd_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 146.000 743.730 154.000 ;
    END
  END s1_wbd_dat_o[22]
  PIN s1_wbd_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 146.000 742.810 154.000 ;
    END
  END s1_wbd_dat_o[23]
  PIN s1_wbd_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 146.000 741.890 154.000 ;
    END
  END s1_wbd_dat_o[24]
  PIN s1_wbd_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 146.000 740.970 154.000 ;
    END
  END s1_wbd_dat_o[25]
  PIN s1_wbd_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 146.000 740.050 154.000 ;
    END
  END s1_wbd_dat_o[26]
  PIN s1_wbd_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.850 146.000 739.130 154.000 ;
    END
  END s1_wbd_dat_o[27]
  PIN s1_wbd_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 146.000 738.210 154.000 ;
    END
  END s1_wbd_dat_o[28]
  PIN s1_wbd_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 146.000 737.290 154.000 ;
    END
  END s1_wbd_dat_o[29]
  PIN s1_wbd_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.850 146.000 762.130 154.000 ;
    END
  END s1_wbd_dat_o[2]
  PIN s1_wbd_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.090 146.000 736.370 154.000 ;
    END
  END s1_wbd_dat_o[30]
  PIN s1_wbd_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 146.000 735.450 154.000 ;
    END
  END s1_wbd_dat_o[31]
  PIN s1_wbd_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930 146.000 761.210 154.000 ;
    END
  END s1_wbd_dat_o[3]
  PIN s1_wbd_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 146.000 760.290 154.000 ;
    END
  END s1_wbd_dat_o[4]
  PIN s1_wbd_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 146.000 759.370 154.000 ;
    END
  END s1_wbd_dat_o[5]
  PIN s1_wbd_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 146.000 758.450 154.000 ;
    END
  END s1_wbd_dat_o[6]
  PIN s1_wbd_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 146.000 757.530 154.000 ;
    END
  END s1_wbd_dat_o[7]
  PIN s1_wbd_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.330 146.000 756.610 154.000 ;
    END
  END s1_wbd_dat_o[8]
  PIN s1_wbd_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.410 146.000 755.690 154.000 ;
    END
  END s1_wbd_dat_o[9]
  PIN s1_wbd_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 146.000 734.530 154.000 ;
    END
  END s1_wbd_sel_o[0]
  PIN s1_wbd_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 146.000 733.610 154.000 ;
    END
  END s1_wbd_sel_o[1]
  PIN s1_wbd_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 146.000 732.690 154.000 ;
    END
  END s1_wbd_sel_o[2]
  PIN s1_wbd_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 146.000 731.770 154.000 ;
    END
  END s1_wbd_sel_o[3]
  PIN s1_wbd_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 146.000 700.490 154.000 ;
    END
  END s1_wbd_stb_o
  PIN s1_wbd_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 146.000 701.410 154.000 ;
    END
  END s1_wbd_we_o
  PIN s2_wbd_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1772.010 146.000 1772.290 154.000 ;
    END
  END s2_wbd_ack_i
  PIN s2_wbd_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1708.530 146.000 1708.810 154.000 ;
    END
  END s2_wbd_adr_o[0]
  PIN s2_wbd_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1707.610 146.000 1707.890 154.000 ;
    END
  END s2_wbd_adr_o[1]
  PIN s2_wbd_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.690 146.000 1706.970 154.000 ;
    END
  END s2_wbd_adr_o[2]
  PIN s2_wbd_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.770 146.000 1706.050 154.000 ;
    END
  END s2_wbd_adr_o[3]
  PIN s2_wbd_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.850 146.000 1705.130 154.000 ;
    END
  END s2_wbd_adr_o[4]
  PIN s2_wbd_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.930 146.000 1704.210 154.000 ;
    END
  END s2_wbd_adr_o[5]
  PIN s2_wbd_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.010 146.000 1703.290 154.000 ;
    END
  END s2_wbd_adr_o[6]
  PIN s2_wbd_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.090 146.000 1702.370 154.000 ;
    END
  END s2_wbd_adr_o[7]
  PIN s2_wbd_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1772.930 146.000 1773.210 154.000 ;
    END
  END s2_wbd_cyc_o
  PIN s2_wbd_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.090 146.000 1771.370 154.000 ;
    END
  END s2_wbd_dat_i[0]
  PIN s2_wbd_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.890 146.000 1762.170 154.000 ;
    END
  END s2_wbd_dat_i[10]
  PIN s2_wbd_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.970 146.000 1761.250 154.000 ;
    END
  END s2_wbd_dat_i[11]
  PIN s2_wbd_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.050 146.000 1760.330 154.000 ;
    END
  END s2_wbd_dat_i[12]
  PIN s2_wbd_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1759.130 146.000 1759.410 154.000 ;
    END
  END s2_wbd_dat_i[13]
  PIN s2_wbd_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.210 146.000 1758.490 154.000 ;
    END
  END s2_wbd_dat_i[14]
  PIN s2_wbd_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1757.290 146.000 1757.570 154.000 ;
    END
  END s2_wbd_dat_i[15]
  PIN s2_wbd_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.370 146.000 1756.650 154.000 ;
    END
  END s2_wbd_dat_i[16]
  PIN s2_wbd_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1755.450 146.000 1755.730 154.000 ;
    END
  END s2_wbd_dat_i[17]
  PIN s2_wbd_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.530 146.000 1754.810 154.000 ;
    END
  END s2_wbd_dat_i[18]
  PIN s2_wbd_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1753.610 146.000 1753.890 154.000 ;
    END
  END s2_wbd_dat_i[19]
  PIN s2_wbd_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.170 146.000 1770.450 154.000 ;
    END
  END s2_wbd_dat_i[1]
  PIN s2_wbd_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.690 146.000 1752.970 154.000 ;
    END
  END s2_wbd_dat_i[20]
  PIN s2_wbd_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.770 146.000 1752.050 154.000 ;
    END
  END s2_wbd_dat_i[21]
  PIN s2_wbd_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1750.850 146.000 1751.130 154.000 ;
    END
  END s2_wbd_dat_i[22]
  PIN s2_wbd_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.930 146.000 1750.210 154.000 ;
    END
  END s2_wbd_dat_i[23]
  PIN s2_wbd_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.010 146.000 1749.290 154.000 ;
    END
  END s2_wbd_dat_i[24]
  PIN s2_wbd_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1748.090 146.000 1748.370 154.000 ;
    END
  END s2_wbd_dat_i[25]
  PIN s2_wbd_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.170 146.000 1747.450 154.000 ;
    END
  END s2_wbd_dat_i[26]
  PIN s2_wbd_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.250 146.000 1746.530 154.000 ;
    END
  END s2_wbd_dat_i[27]
  PIN s2_wbd_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.330 146.000 1745.610 154.000 ;
    END
  END s2_wbd_dat_i[28]
  PIN s2_wbd_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1744.410 146.000 1744.690 154.000 ;
    END
  END s2_wbd_dat_i[29]
  PIN s2_wbd_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1769.250 146.000 1769.530 154.000 ;
    END
  END s2_wbd_dat_i[2]
  PIN s2_wbd_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.490 146.000 1743.770 154.000 ;
    END
  END s2_wbd_dat_i[30]
  PIN s2_wbd_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.570 146.000 1742.850 154.000 ;
    END
  END s2_wbd_dat_i[31]
  PIN s2_wbd_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1768.330 146.000 1768.610 154.000 ;
    END
  END s2_wbd_dat_i[3]
  PIN s2_wbd_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1767.410 146.000 1767.690 154.000 ;
    END
  END s2_wbd_dat_i[4]
  PIN s2_wbd_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1766.490 146.000 1766.770 154.000 ;
    END
  END s2_wbd_dat_i[5]
  PIN s2_wbd_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.570 146.000 1765.850 154.000 ;
    END
  END s2_wbd_dat_i[6]
  PIN s2_wbd_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.650 146.000 1764.930 154.000 ;
    END
  END s2_wbd_dat_i[7]
  PIN s2_wbd_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1763.730 146.000 1764.010 154.000 ;
    END
  END s2_wbd_dat_i[8]
  PIN s2_wbd_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.810 146.000 1763.090 154.000 ;
    END
  END s2_wbd_dat_i[9]
  PIN s2_wbd_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1741.650 146.000 1741.930 154.000 ;
    END
  END s2_wbd_dat_o[0]
  PIN s2_wbd_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.450 146.000 1732.730 154.000 ;
    END
  END s2_wbd_dat_o[10]
  PIN s2_wbd_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1731.530 146.000 1731.810 154.000 ;
    END
  END s2_wbd_dat_o[11]
  PIN s2_wbd_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1730.610 146.000 1730.890 154.000 ;
    END
  END s2_wbd_dat_o[12]
  PIN s2_wbd_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.690 146.000 1729.970 154.000 ;
    END
  END s2_wbd_dat_o[13]
  PIN s2_wbd_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.770 146.000 1729.050 154.000 ;
    END
  END s2_wbd_dat_o[14]
  PIN s2_wbd_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.850 146.000 1728.130 154.000 ;
    END
  END s2_wbd_dat_o[15]
  PIN s2_wbd_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.930 146.000 1727.210 154.000 ;
    END
  END s2_wbd_dat_o[16]
  PIN s2_wbd_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.010 146.000 1726.290 154.000 ;
    END
  END s2_wbd_dat_o[17]
  PIN s2_wbd_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1725.090 146.000 1725.370 154.000 ;
    END
  END s2_wbd_dat_o[18]
  PIN s2_wbd_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1724.170 146.000 1724.450 154.000 ;
    END
  END s2_wbd_dat_o[19]
  PIN s2_wbd_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.730 146.000 1741.010 154.000 ;
    END
  END s2_wbd_dat_o[1]
  PIN s2_wbd_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1723.250 146.000 1723.530 154.000 ;
    END
  END s2_wbd_dat_o[20]
  PIN s2_wbd_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.330 146.000 1722.610 154.000 ;
    END
  END s2_wbd_dat_o[21]
  PIN s2_wbd_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.410 146.000 1721.690 154.000 ;
    END
  END s2_wbd_dat_o[22]
  PIN s2_wbd_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1720.490 146.000 1720.770 154.000 ;
    END
  END s2_wbd_dat_o[23]
  PIN s2_wbd_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.570 146.000 1719.850 154.000 ;
    END
  END s2_wbd_dat_o[24]
  PIN s2_wbd_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.650 146.000 1718.930 154.000 ;
    END
  END s2_wbd_dat_o[25]
  PIN s2_wbd_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1717.730 146.000 1718.010 154.000 ;
    END
  END s2_wbd_dat_o[26]
  PIN s2_wbd_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.810 146.000 1717.090 154.000 ;
    END
  END s2_wbd_dat_o[27]
  PIN s2_wbd_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.890 146.000 1716.170 154.000 ;
    END
  END s2_wbd_dat_o[28]
  PIN s2_wbd_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.970 146.000 1715.250 154.000 ;
    END
  END s2_wbd_dat_o[29]
  PIN s2_wbd_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.810 146.000 1740.090 154.000 ;
    END
  END s2_wbd_dat_o[2]
  PIN s2_wbd_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.050 146.000 1714.330 154.000 ;
    END
  END s2_wbd_dat_o[30]
  PIN s2_wbd_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.130 146.000 1713.410 154.000 ;
    END
  END s2_wbd_dat_o[31]
  PIN s2_wbd_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.890 146.000 1739.170 154.000 ;
    END
  END s2_wbd_dat_o[3]
  PIN s2_wbd_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.970 146.000 1738.250 154.000 ;
    END
  END s2_wbd_dat_o[4]
  PIN s2_wbd_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.050 146.000 1737.330 154.000 ;
    END
  END s2_wbd_dat_o[5]
  PIN s2_wbd_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.130 146.000 1736.410 154.000 ;
    END
  END s2_wbd_dat_o[6]
  PIN s2_wbd_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.210 146.000 1735.490 154.000 ;
    END
  END s2_wbd_dat_o[7]
  PIN s2_wbd_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.290 146.000 1734.570 154.000 ;
    END
  END s2_wbd_dat_o[8]
  PIN s2_wbd_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.370 146.000 1733.650 154.000 ;
    END
  END s2_wbd_dat_o[9]
  PIN s2_wbd_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.210 146.000 1712.490 154.000 ;
    END
  END s2_wbd_sel_o[0]
  PIN s2_wbd_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.290 146.000 1711.570 154.000 ;
    END
  END s2_wbd_sel_o[1]
  PIN s2_wbd_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.370 146.000 1710.650 154.000 ;
    END
  END s2_wbd_sel_o[2]
  PIN s2_wbd_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.450 146.000 1709.730 154.000 ;
    END
  END s2_wbd_sel_o[3]
  PIN s2_wbd_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 146.000 1700.530 154.000 ;
    END
  END s2_wbd_stb_o
  PIN s2_wbd_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1701.170 146.000 1701.450 154.000 ;
    END
  END s2_wbd_we_o
  PIN s3_wbd_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.110 -4.000 1972.390 4.000 ;
    END
  END s3_wbd_ack_i
  PIN s3_wbd_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1908.630 -4.000 1908.910 4.000 ;
    END
  END s3_wbd_adr_o[0]
  PIN s3_wbd_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1907.710 -4.000 1907.990 4.000 ;
    END
  END s3_wbd_adr_o[1]
  PIN s3_wbd_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1906.790 -4.000 1907.070 4.000 ;
    END
  END s3_wbd_adr_o[2]
  PIN s3_wbd_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.870 -4.000 1906.150 4.000 ;
    END
  END s3_wbd_adr_o[3]
  PIN s3_wbd_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.950 -4.000 1905.230 4.000 ;
    END
  END s3_wbd_adr_o[4]
  PIN s3_wbd_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.030 -4.000 1904.310 4.000 ;
    END
  END s3_wbd_adr_o[5]
  PIN s3_wbd_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.110 -4.000 1903.390 4.000 ;
    END
  END s3_wbd_adr_o[6]
  PIN s3_wbd_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1902.190 -4.000 1902.470 4.000 ;
    END
  END s3_wbd_adr_o[7]
  PIN s3_wbd_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1973.030 -4.000 1973.310 4.000 ;
    END
  END s3_wbd_cyc_o
  PIN s3_wbd_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.190 -4.000 1971.470 4.000 ;
    END
  END s3_wbd_dat_i[0]
  PIN s3_wbd_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.990 -4.000 1962.270 4.000 ;
    END
  END s3_wbd_dat_i[10]
  PIN s3_wbd_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.070 -4.000 1961.350 4.000 ;
    END
  END s3_wbd_dat_i[11]
  PIN s3_wbd_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1960.150 -4.000 1960.430 4.000 ;
    END
  END s3_wbd_dat_i[12]
  PIN s3_wbd_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.230 -4.000 1959.510 4.000 ;
    END
  END s3_wbd_dat_i[13]
  PIN s3_wbd_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1958.310 -4.000 1958.590 4.000 ;
    END
  END s3_wbd_dat_i[14]
  PIN s3_wbd_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1957.390 -4.000 1957.670 4.000 ;
    END
  END s3_wbd_dat_i[15]
  PIN s3_wbd_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.470 -4.000 1956.750 4.000 ;
    END
  END s3_wbd_dat_i[16]
  PIN s3_wbd_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1955.550 -4.000 1955.830 4.000 ;
    END
  END s3_wbd_dat_i[17]
  PIN s3_wbd_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.630 -4.000 1954.910 4.000 ;
    END
  END s3_wbd_dat_i[18]
  PIN s3_wbd_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.710 -4.000 1953.990 4.000 ;
    END
  END s3_wbd_dat_i[19]
  PIN s3_wbd_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1970.270 -4.000 1970.550 4.000 ;
    END
  END s3_wbd_dat_i[1]
  PIN s3_wbd_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1952.790 -4.000 1953.070 4.000 ;
    END
  END s3_wbd_dat_i[20]
  PIN s3_wbd_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1951.870 -4.000 1952.150 4.000 ;
    END
  END s3_wbd_dat_i[21]
  PIN s3_wbd_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1950.950 -4.000 1951.230 4.000 ;
    END
  END s3_wbd_dat_i[22]
  PIN s3_wbd_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1950.030 -4.000 1950.310 4.000 ;
    END
  END s3_wbd_dat_i[23]
  PIN s3_wbd_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1949.110 -4.000 1949.390 4.000 ;
    END
  END s3_wbd_dat_i[24]
  PIN s3_wbd_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.190 -4.000 1948.470 4.000 ;
    END
  END s3_wbd_dat_i[25]
  PIN s3_wbd_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.270 -4.000 1947.550 4.000 ;
    END
  END s3_wbd_dat_i[26]
  PIN s3_wbd_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1946.350 -4.000 1946.630 4.000 ;
    END
  END s3_wbd_dat_i[27]
  PIN s3_wbd_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.430 -4.000 1945.710 4.000 ;
    END
  END s3_wbd_dat_i[28]
  PIN s3_wbd_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1944.510 -4.000 1944.790 4.000 ;
    END
  END s3_wbd_dat_i[29]
  PIN s3_wbd_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1969.350 -4.000 1969.630 4.000 ;
    END
  END s3_wbd_dat_i[2]
  PIN s3_wbd_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1943.590 -4.000 1943.870 4.000 ;
    END
  END s3_wbd_dat_i[30]
  PIN s3_wbd_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1942.670 -4.000 1942.950 4.000 ;
    END
  END s3_wbd_dat_i[31]
  PIN s3_wbd_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1968.430 -4.000 1968.710 4.000 ;
    END
  END s3_wbd_dat_i[3]
  PIN s3_wbd_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.510 -4.000 1967.790 4.000 ;
    END
  END s3_wbd_dat_i[4]
  PIN s3_wbd_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1966.590 -4.000 1966.870 4.000 ;
    END
  END s3_wbd_dat_i[5]
  PIN s3_wbd_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.670 -4.000 1965.950 4.000 ;
    END
  END s3_wbd_dat_i[6]
  PIN s3_wbd_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1964.750 -4.000 1965.030 4.000 ;
    END
  END s3_wbd_dat_i[7]
  PIN s3_wbd_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1963.830 -4.000 1964.110 4.000 ;
    END
  END s3_wbd_dat_i[8]
  PIN s3_wbd_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1962.910 -4.000 1963.190 4.000 ;
    END
  END s3_wbd_dat_i[9]
  PIN s3_wbd_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.750 -4.000 1942.030 4.000 ;
    END
  END s3_wbd_dat_o[0]
  PIN s3_wbd_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.550 -4.000 1932.830 4.000 ;
    END
  END s3_wbd_dat_o[10]
  PIN s3_wbd_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1931.630 -4.000 1931.910 4.000 ;
    END
  END s3_wbd_dat_o[11]
  PIN s3_wbd_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1930.710 -4.000 1930.990 4.000 ;
    END
  END s3_wbd_dat_o[12]
  PIN s3_wbd_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.790 -4.000 1930.070 4.000 ;
    END
  END s3_wbd_dat_o[13]
  PIN s3_wbd_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1928.870 -4.000 1929.150 4.000 ;
    END
  END s3_wbd_dat_o[14]
  PIN s3_wbd_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.950 -4.000 1928.230 4.000 ;
    END
  END s3_wbd_dat_o[15]
  PIN s3_wbd_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.030 -4.000 1927.310 4.000 ;
    END
  END s3_wbd_dat_o[16]
  PIN s3_wbd_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1926.110 -4.000 1926.390 4.000 ;
    END
  END s3_wbd_dat_o[17]
  PIN s3_wbd_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1925.190 -4.000 1925.470 4.000 ;
    END
  END s3_wbd_dat_o[18]
  PIN s3_wbd_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1924.270 -4.000 1924.550 4.000 ;
    END
  END s3_wbd_dat_o[19]
  PIN s3_wbd_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1940.830 -4.000 1941.110 4.000 ;
    END
  END s3_wbd_dat_o[1]
  PIN s3_wbd_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.350 -4.000 1923.630 4.000 ;
    END
  END s3_wbd_dat_o[20]
  PIN s3_wbd_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.430 -4.000 1922.710 4.000 ;
    END
  END s3_wbd_dat_o[21]
  PIN s3_wbd_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1921.510 -4.000 1921.790 4.000 ;
    END
  END s3_wbd_dat_o[22]
  PIN s3_wbd_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1920.590 -4.000 1920.870 4.000 ;
    END
  END s3_wbd_dat_o[23]
  PIN s3_wbd_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.670 -4.000 1919.950 4.000 ;
    END
  END s3_wbd_dat_o[24]
  PIN s3_wbd_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1918.750 -4.000 1919.030 4.000 ;
    END
  END s3_wbd_dat_o[25]
  PIN s3_wbd_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.830 -4.000 1918.110 4.000 ;
    END
  END s3_wbd_dat_o[26]
  PIN s3_wbd_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1916.910 -4.000 1917.190 4.000 ;
    END
  END s3_wbd_dat_o[27]
  PIN s3_wbd_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.990 -4.000 1916.270 4.000 ;
    END
  END s3_wbd_dat_o[28]
  PIN s3_wbd_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.070 -4.000 1915.350 4.000 ;
    END
  END s3_wbd_dat_o[29]
  PIN s3_wbd_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1939.910 -4.000 1940.190 4.000 ;
    END
  END s3_wbd_dat_o[2]
  PIN s3_wbd_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1914.150 -4.000 1914.430 4.000 ;
    END
  END s3_wbd_dat_o[30]
  PIN s3_wbd_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1913.230 -4.000 1913.510 4.000 ;
    END
  END s3_wbd_dat_o[31]
  PIN s3_wbd_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.990 -4.000 1939.270 4.000 ;
    END
  END s3_wbd_dat_o[3]
  PIN s3_wbd_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.070 -4.000 1938.350 4.000 ;
    END
  END s3_wbd_dat_o[4]
  PIN s3_wbd_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1937.150 -4.000 1937.430 4.000 ;
    END
  END s3_wbd_dat_o[5]
  PIN s3_wbd_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1936.230 -4.000 1936.510 4.000 ;
    END
  END s3_wbd_dat_o[6]
  PIN s3_wbd_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.310 -4.000 1935.590 4.000 ;
    END
  END s3_wbd_dat_o[7]
  PIN s3_wbd_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1934.390 -4.000 1934.670 4.000 ;
    END
  END s3_wbd_dat_o[8]
  PIN s3_wbd_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.470 -4.000 1933.750 4.000 ;
    END
  END s3_wbd_dat_o[9]
  PIN s3_wbd_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.310 -4.000 1912.590 4.000 ;
    END
  END s3_wbd_sel_o[0]
  PIN s3_wbd_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.390 -4.000 1911.670 4.000 ;
    END
  END s3_wbd_sel_o[1]
  PIN s3_wbd_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1910.470 -4.000 1910.750 4.000 ;
    END
  END s3_wbd_sel_o[2]
  PIN s3_wbd_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.550 -4.000 1909.830 4.000 ;
    END
  END s3_wbd_sel_o[3]
  PIN s3_wbd_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1900.350 -4.000 1900.630 4.000 ;
    END
  END s3_wbd_stb_o
  PIN s3_wbd_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1901.270 -4.000 1901.550 4.000 ;
    END
  END s3_wbd_we_o
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1828.155 10.640 1831.155 138.960 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1098.500 10.640 1101.500 138.960 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 368.845 10.640 371.845 138.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1463.325 10.640 1466.325 138.960 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 733.675 10.640 736.675 138.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 0.425 2194.200 149.515 ;
      LAYER met1 ;
        RECT 0.530 0.040 2194.200 149.560 ;
      LAYER met2 ;
        RECT 1.110 145.720 1.190 149.590 ;
        RECT 2.030 145.720 2.110 149.590 ;
        RECT 2.950 145.720 3.030 149.590 ;
        RECT 3.870 145.720 3.950 149.590 ;
        RECT 4.790 145.720 4.870 149.590 ;
        RECT 5.710 145.720 5.790 149.590 ;
        RECT 6.630 145.720 6.710 149.590 ;
        RECT 7.550 145.720 7.630 149.590 ;
        RECT 8.470 145.720 8.550 149.590 ;
        RECT 9.390 145.720 9.470 149.590 ;
        RECT 10.310 145.720 10.390 149.590 ;
        RECT 11.230 145.720 11.310 149.590 ;
        RECT 12.150 145.720 12.230 149.590 ;
        RECT 13.070 145.720 13.150 149.590 ;
        RECT 13.990 145.720 14.070 149.590 ;
        RECT 14.910 145.720 14.990 149.590 ;
        RECT 15.830 145.720 15.910 149.590 ;
        RECT 16.750 145.720 16.830 149.590 ;
        RECT 17.670 145.720 17.750 149.590 ;
        RECT 18.590 145.720 18.670 149.590 ;
        RECT 19.510 145.720 19.590 149.590 ;
        RECT 20.430 145.720 20.510 149.590 ;
        RECT 21.350 145.720 21.430 149.590 ;
        RECT 22.270 145.720 22.350 149.590 ;
        RECT 23.190 145.720 23.270 149.590 ;
        RECT 24.110 145.720 24.190 149.590 ;
        RECT 25.030 145.720 25.110 149.590 ;
        RECT 25.950 145.720 26.030 149.590 ;
        RECT 26.870 145.720 26.950 149.590 ;
        RECT 27.790 145.720 27.870 149.590 ;
        RECT 28.710 145.720 28.790 149.590 ;
        RECT 29.630 145.720 29.710 149.590 ;
        RECT 30.550 145.720 30.630 149.590 ;
        RECT 31.470 145.720 31.550 149.590 ;
        RECT 32.390 145.720 32.470 149.590 ;
        RECT 33.310 145.720 33.390 149.590 ;
        RECT 34.230 145.720 34.310 149.590 ;
        RECT 35.150 145.720 35.230 149.590 ;
        RECT 36.070 145.720 36.150 149.590 ;
        RECT 36.990 145.720 37.070 149.590 ;
        RECT 37.910 145.720 37.990 149.590 ;
        RECT 38.830 145.720 38.910 149.590 ;
        RECT 39.750 145.720 39.830 149.590 ;
        RECT 40.670 145.720 40.750 149.590 ;
        RECT 41.590 145.720 41.670 149.590 ;
        RECT 42.510 145.720 42.590 149.590 ;
        RECT 43.430 145.720 43.510 149.590 ;
        RECT 44.350 145.720 44.430 149.590 ;
        RECT 45.270 145.720 45.350 149.590 ;
        RECT 46.190 145.720 46.270 149.590 ;
        RECT 47.110 145.720 47.190 149.590 ;
        RECT 48.030 145.720 48.110 149.590 ;
        RECT 48.950 145.720 49.030 149.590 ;
        RECT 49.870 145.720 49.950 149.590 ;
        RECT 50.790 145.720 50.870 149.590 ;
        RECT 51.710 145.720 51.790 149.590 ;
        RECT 52.630 145.720 52.710 149.590 ;
        RECT 53.550 145.720 53.630 149.590 ;
        RECT 54.470 145.720 54.550 149.590 ;
        RECT 55.390 145.720 55.470 149.590 ;
        RECT 56.310 145.720 56.390 149.590 ;
        RECT 57.230 145.720 57.310 149.590 ;
        RECT 58.150 145.720 58.230 149.590 ;
        RECT 59.070 145.720 59.150 149.590 ;
        RECT 59.990 145.720 60.070 149.590 ;
        RECT 60.910 145.720 60.990 149.590 ;
        RECT 61.830 145.720 61.910 149.590 ;
        RECT 62.750 145.720 62.830 149.590 ;
        RECT 63.670 145.720 63.750 149.590 ;
        RECT 64.590 145.720 64.670 149.590 ;
        RECT 65.510 145.720 65.590 149.590 ;
        RECT 66.430 145.720 66.510 149.590 ;
        RECT 67.350 145.720 67.430 149.590 ;
        RECT 68.270 145.720 68.350 149.590 ;
        RECT 69.190 145.720 69.270 149.590 ;
        RECT 70.110 145.720 70.190 149.590 ;
        RECT 71.030 145.720 71.110 149.590 ;
        RECT 71.950 145.720 72.030 149.590 ;
        RECT 72.870 145.720 72.950 149.590 ;
        RECT 73.790 145.720 73.870 149.590 ;
        RECT 74.710 145.720 74.790 149.590 ;
        RECT 75.630 145.720 75.710 149.590 ;
        RECT 76.550 145.720 76.630 149.590 ;
        RECT 77.470 145.720 77.550 149.590 ;
        RECT 78.390 145.720 78.470 149.590 ;
        RECT 79.310 145.720 79.390 149.590 ;
        RECT 80.230 145.720 80.310 149.590 ;
        RECT 81.150 145.720 81.230 149.590 ;
        RECT 82.070 145.720 82.150 149.590 ;
        RECT 82.990 145.720 83.070 149.590 ;
        RECT 83.910 145.720 83.990 149.590 ;
        RECT 84.830 145.720 84.910 149.590 ;
        RECT 85.750 145.720 85.830 149.590 ;
        RECT 86.670 145.720 86.750 149.590 ;
        RECT 87.590 145.720 87.670 149.590 ;
        RECT 88.510 145.720 88.590 149.590 ;
        RECT 89.430 145.720 89.510 149.590 ;
        RECT 90.350 145.720 90.430 149.590 ;
        RECT 91.270 145.720 91.350 149.590 ;
        RECT 92.190 145.720 92.270 149.590 ;
        RECT 93.110 145.720 93.190 149.590 ;
        RECT 94.030 145.720 94.110 149.590 ;
        RECT 94.950 145.720 95.030 149.590 ;
        RECT 95.870 145.720 699.930 149.590 ;
        RECT 700.770 145.720 700.850 149.590 ;
        RECT 701.690 145.720 701.770 149.590 ;
        RECT 702.610 145.720 702.690 149.590 ;
        RECT 703.530 145.720 703.610 149.590 ;
        RECT 704.450 145.720 704.530 149.590 ;
        RECT 705.370 145.720 705.450 149.590 ;
        RECT 706.290 145.720 706.370 149.590 ;
        RECT 707.210 145.720 707.290 149.590 ;
        RECT 708.130 145.720 708.210 149.590 ;
        RECT 709.050 145.720 709.130 149.590 ;
        RECT 709.970 145.720 710.050 149.590 ;
        RECT 710.890 145.720 710.970 149.590 ;
        RECT 711.810 145.720 711.890 149.590 ;
        RECT 712.730 145.720 712.810 149.590 ;
        RECT 713.650 145.720 713.730 149.590 ;
        RECT 714.570 145.720 714.650 149.590 ;
        RECT 715.490 145.720 715.570 149.590 ;
        RECT 716.410 145.720 716.490 149.590 ;
        RECT 717.330 145.720 717.410 149.590 ;
        RECT 718.250 145.720 718.330 149.590 ;
        RECT 719.170 145.720 719.250 149.590 ;
        RECT 720.090 145.720 720.170 149.590 ;
        RECT 721.010 145.720 721.090 149.590 ;
        RECT 721.930 145.720 722.010 149.590 ;
        RECT 722.850 145.720 722.930 149.590 ;
        RECT 723.770 145.720 723.850 149.590 ;
        RECT 724.690 145.720 724.770 149.590 ;
        RECT 725.610 145.720 725.690 149.590 ;
        RECT 726.530 145.720 726.610 149.590 ;
        RECT 727.450 145.720 727.530 149.590 ;
        RECT 728.370 145.720 728.450 149.590 ;
        RECT 729.290 145.720 729.370 149.590 ;
        RECT 730.210 145.720 730.290 149.590 ;
        RECT 731.130 145.720 731.210 149.590 ;
        RECT 732.050 145.720 732.130 149.590 ;
        RECT 732.970 145.720 733.050 149.590 ;
        RECT 733.890 145.720 733.970 149.590 ;
        RECT 734.810 145.720 734.890 149.590 ;
        RECT 735.730 145.720 735.810 149.590 ;
        RECT 736.650 145.720 736.730 149.590 ;
        RECT 737.570 145.720 737.650 149.590 ;
        RECT 738.490 145.720 738.570 149.590 ;
        RECT 739.410 145.720 739.490 149.590 ;
        RECT 740.330 145.720 740.410 149.590 ;
        RECT 741.250 145.720 741.330 149.590 ;
        RECT 742.170 145.720 742.250 149.590 ;
        RECT 743.090 145.720 743.170 149.590 ;
        RECT 744.010 145.720 744.090 149.590 ;
        RECT 744.930 145.720 745.010 149.590 ;
        RECT 745.850 145.720 745.930 149.590 ;
        RECT 746.770 145.720 746.850 149.590 ;
        RECT 747.690 145.720 747.770 149.590 ;
        RECT 748.610 145.720 748.690 149.590 ;
        RECT 749.530 145.720 749.610 149.590 ;
        RECT 750.450 145.720 750.530 149.590 ;
        RECT 751.370 145.720 751.450 149.590 ;
        RECT 752.290 145.720 752.370 149.590 ;
        RECT 753.210 145.720 753.290 149.590 ;
        RECT 754.130 145.720 754.210 149.590 ;
        RECT 755.050 145.720 755.130 149.590 ;
        RECT 755.970 145.720 756.050 149.590 ;
        RECT 756.890 145.720 756.970 149.590 ;
        RECT 757.810 145.720 757.890 149.590 ;
        RECT 758.730 145.720 758.810 149.590 ;
        RECT 759.650 145.720 759.730 149.590 ;
        RECT 760.570 145.720 760.650 149.590 ;
        RECT 761.490 145.720 761.570 149.590 ;
        RECT 762.410 145.720 762.490 149.590 ;
        RECT 763.330 145.720 763.410 149.590 ;
        RECT 764.250 145.720 764.330 149.590 ;
        RECT 765.170 145.720 765.250 149.590 ;
        RECT 766.090 145.720 766.170 149.590 ;
        RECT 767.010 145.720 767.090 149.590 ;
        RECT 767.930 145.720 768.010 149.590 ;
        RECT 768.850 145.720 768.930 149.590 ;
        RECT 769.770 145.720 769.850 149.590 ;
        RECT 770.690 145.720 770.770 149.590 ;
        RECT 771.610 145.720 771.690 149.590 ;
        RECT 772.530 145.720 772.610 149.590 ;
        RECT 773.450 145.720 773.530 149.590 ;
        RECT 774.370 145.720 774.450 149.590 ;
        RECT 775.290 145.720 775.370 149.590 ;
        RECT 776.210 145.720 776.290 149.590 ;
        RECT 777.130 145.720 777.210 149.590 ;
        RECT 778.050 145.720 778.130 149.590 ;
        RECT 778.970 145.720 779.050 149.590 ;
        RECT 779.890 145.720 779.970 149.590 ;
        RECT 780.810 145.720 780.890 149.590 ;
        RECT 781.730 145.720 781.810 149.590 ;
        RECT 782.650 145.720 782.730 149.590 ;
        RECT 783.570 145.720 783.650 149.590 ;
        RECT 784.490 145.720 784.570 149.590 ;
        RECT 785.410 145.720 785.490 149.590 ;
        RECT 786.330 145.720 786.410 149.590 ;
        RECT 787.250 145.720 787.330 149.590 ;
        RECT 788.170 145.720 788.250 149.590 ;
        RECT 789.090 145.720 789.170 149.590 ;
        RECT 790.010 145.720 790.090 149.590 ;
        RECT 790.930 145.720 791.010 149.590 ;
        RECT 791.850 145.720 791.930 149.590 ;
        RECT 792.770 145.720 792.850 149.590 ;
        RECT 793.690 145.720 793.770 149.590 ;
        RECT 794.610 145.720 794.690 149.590 ;
        RECT 795.530 145.720 1699.970 149.590 ;
        RECT 1700.810 145.720 1700.890 149.590 ;
        RECT 1701.730 145.720 1701.810 149.590 ;
        RECT 1702.650 145.720 1702.730 149.590 ;
        RECT 1703.570 145.720 1703.650 149.590 ;
        RECT 1704.490 145.720 1704.570 149.590 ;
        RECT 1705.410 145.720 1705.490 149.590 ;
        RECT 1706.330 145.720 1706.410 149.590 ;
        RECT 1707.250 145.720 1707.330 149.590 ;
        RECT 1708.170 145.720 1708.250 149.590 ;
        RECT 1709.090 145.720 1709.170 149.590 ;
        RECT 1710.010 145.720 1710.090 149.590 ;
        RECT 1710.930 145.720 1711.010 149.590 ;
        RECT 1711.850 145.720 1711.930 149.590 ;
        RECT 1712.770 145.720 1712.850 149.590 ;
        RECT 1713.690 145.720 1713.770 149.590 ;
        RECT 1714.610 145.720 1714.690 149.590 ;
        RECT 1715.530 145.720 1715.610 149.590 ;
        RECT 1716.450 145.720 1716.530 149.590 ;
        RECT 1717.370 145.720 1717.450 149.590 ;
        RECT 1718.290 145.720 1718.370 149.590 ;
        RECT 1719.210 145.720 1719.290 149.590 ;
        RECT 1720.130 145.720 1720.210 149.590 ;
        RECT 1721.050 145.720 1721.130 149.590 ;
        RECT 1721.970 145.720 1722.050 149.590 ;
        RECT 1722.890 145.720 1722.970 149.590 ;
        RECT 1723.810 145.720 1723.890 149.590 ;
        RECT 1724.730 145.720 1724.810 149.590 ;
        RECT 1725.650 145.720 1725.730 149.590 ;
        RECT 1726.570 145.720 1726.650 149.590 ;
        RECT 1727.490 145.720 1727.570 149.590 ;
        RECT 1728.410 145.720 1728.490 149.590 ;
        RECT 1729.330 145.720 1729.410 149.590 ;
        RECT 1730.250 145.720 1730.330 149.590 ;
        RECT 1731.170 145.720 1731.250 149.590 ;
        RECT 1732.090 145.720 1732.170 149.590 ;
        RECT 1733.010 145.720 1733.090 149.590 ;
        RECT 1733.930 145.720 1734.010 149.590 ;
        RECT 1734.850 145.720 1734.930 149.590 ;
        RECT 1735.770 145.720 1735.850 149.590 ;
        RECT 1736.690 145.720 1736.770 149.590 ;
        RECT 1737.610 145.720 1737.690 149.590 ;
        RECT 1738.530 145.720 1738.610 149.590 ;
        RECT 1739.450 145.720 1739.530 149.590 ;
        RECT 1740.370 145.720 1740.450 149.590 ;
        RECT 1741.290 145.720 1741.370 149.590 ;
        RECT 1742.210 145.720 1742.290 149.590 ;
        RECT 1743.130 145.720 1743.210 149.590 ;
        RECT 1744.050 145.720 1744.130 149.590 ;
        RECT 1744.970 145.720 1745.050 149.590 ;
        RECT 1745.890 145.720 1745.970 149.590 ;
        RECT 1746.810 145.720 1746.890 149.590 ;
        RECT 1747.730 145.720 1747.810 149.590 ;
        RECT 1748.650 145.720 1748.730 149.590 ;
        RECT 1749.570 145.720 1749.650 149.590 ;
        RECT 1750.490 145.720 1750.570 149.590 ;
        RECT 1751.410 145.720 1751.490 149.590 ;
        RECT 1752.330 145.720 1752.410 149.590 ;
        RECT 1753.250 145.720 1753.330 149.590 ;
        RECT 1754.170 145.720 1754.250 149.590 ;
        RECT 1755.090 145.720 1755.170 149.590 ;
        RECT 1756.010 145.720 1756.090 149.590 ;
        RECT 1756.930 145.720 1757.010 149.590 ;
        RECT 1757.850 145.720 1757.930 149.590 ;
        RECT 1758.770 145.720 1758.850 149.590 ;
        RECT 1759.690 145.720 1759.770 149.590 ;
        RECT 1760.610 145.720 1760.690 149.590 ;
        RECT 1761.530 145.720 1761.610 149.590 ;
        RECT 1762.450 145.720 1762.530 149.590 ;
        RECT 1763.370 145.720 1763.450 149.590 ;
        RECT 1764.290 145.720 1764.370 149.590 ;
        RECT 1765.210 145.720 1765.290 149.590 ;
        RECT 1766.130 145.720 1766.210 149.590 ;
        RECT 1767.050 145.720 1767.130 149.590 ;
        RECT 1767.970 145.720 1768.050 149.590 ;
        RECT 1768.890 145.720 1768.970 149.590 ;
        RECT 1769.810 145.720 1769.890 149.590 ;
        RECT 1770.730 145.720 1770.810 149.590 ;
        RECT 1771.650 145.720 1771.730 149.590 ;
        RECT 1772.570 145.720 1772.650 149.590 ;
        RECT 1773.490 145.720 2178.010 149.590 ;
        RECT 0.550 4.280 2178.010 145.720 ;
        RECT 1.110 0.010 1.190 4.280 ;
        RECT 2.030 0.010 2.110 4.280 ;
        RECT 2.950 0.010 3.030 4.280 ;
        RECT 3.870 0.010 3.950 4.280 ;
        RECT 4.790 0.010 4.870 4.280 ;
        RECT 5.710 0.010 5.790 4.280 ;
        RECT 6.630 0.010 6.710 4.280 ;
        RECT 7.550 0.010 7.630 4.280 ;
        RECT 8.470 0.010 8.550 4.280 ;
        RECT 9.390 0.010 9.470 4.280 ;
        RECT 10.310 0.010 10.390 4.280 ;
        RECT 11.230 0.010 11.310 4.280 ;
        RECT 12.150 0.010 12.230 4.280 ;
        RECT 13.070 0.010 13.150 4.280 ;
        RECT 13.990 0.010 14.070 4.280 ;
        RECT 14.910 0.010 14.990 4.280 ;
        RECT 15.830 0.010 15.910 4.280 ;
        RECT 16.750 0.010 16.830 4.280 ;
        RECT 17.670 0.010 17.750 4.280 ;
        RECT 18.590 0.010 18.670 4.280 ;
        RECT 19.510 0.010 19.590 4.280 ;
        RECT 20.430 0.010 20.510 4.280 ;
        RECT 21.350 0.010 21.430 4.280 ;
        RECT 22.270 0.010 22.350 4.280 ;
        RECT 23.190 0.010 23.270 4.280 ;
        RECT 24.110 0.010 24.190 4.280 ;
        RECT 25.030 0.010 25.110 4.280 ;
        RECT 25.950 0.010 26.030 4.280 ;
        RECT 26.870 0.010 26.950 4.280 ;
        RECT 27.790 0.010 27.870 4.280 ;
        RECT 28.710 0.010 28.790 4.280 ;
        RECT 29.630 0.010 29.710 4.280 ;
        RECT 30.550 0.010 30.630 4.280 ;
        RECT 31.470 0.010 31.550 4.280 ;
        RECT 32.390 0.010 32.470 4.280 ;
        RECT 33.310 0.010 33.390 4.280 ;
        RECT 34.230 0.010 34.310 4.280 ;
        RECT 35.150 0.010 35.230 4.280 ;
        RECT 36.070 0.010 36.150 4.280 ;
        RECT 36.990 0.010 37.070 4.280 ;
        RECT 37.910 0.010 37.990 4.280 ;
        RECT 38.830 0.010 38.910 4.280 ;
        RECT 39.750 0.010 39.830 4.280 ;
        RECT 40.670 0.010 40.750 4.280 ;
        RECT 41.590 0.010 41.670 4.280 ;
        RECT 42.510 0.010 42.590 4.280 ;
        RECT 43.430 0.010 43.510 4.280 ;
        RECT 44.350 0.010 44.430 4.280 ;
        RECT 45.270 0.010 45.350 4.280 ;
        RECT 46.190 0.010 46.270 4.280 ;
        RECT 47.110 0.010 47.190 4.280 ;
        RECT 48.030 0.010 48.110 4.280 ;
        RECT 48.950 0.010 49.030 4.280 ;
        RECT 49.870 0.010 49.950 4.280 ;
        RECT 50.790 0.010 50.870 4.280 ;
        RECT 51.710 0.010 51.790 4.280 ;
        RECT 52.630 0.010 52.710 4.280 ;
        RECT 53.550 0.010 53.630 4.280 ;
        RECT 54.470 0.010 54.550 4.280 ;
        RECT 55.390 0.010 55.470 4.280 ;
        RECT 56.310 0.010 56.390 4.280 ;
        RECT 57.230 0.010 57.310 4.280 ;
        RECT 58.150 0.010 58.230 4.280 ;
        RECT 59.070 0.010 59.150 4.280 ;
        RECT 59.990 0.010 60.070 4.280 ;
        RECT 60.910 0.010 60.990 4.280 ;
        RECT 61.830 0.010 61.910 4.280 ;
        RECT 62.750 0.010 62.830 4.280 ;
        RECT 63.670 0.010 63.750 4.280 ;
        RECT 64.590 0.010 64.670 4.280 ;
        RECT 65.510 0.010 65.590 4.280 ;
        RECT 66.430 0.010 66.510 4.280 ;
        RECT 67.350 0.010 67.430 4.280 ;
        RECT 68.270 0.010 68.350 4.280 ;
        RECT 69.190 0.010 69.270 4.280 ;
        RECT 70.110 0.010 70.190 4.280 ;
        RECT 71.030 0.010 71.110 4.280 ;
        RECT 71.950 0.010 72.030 4.280 ;
        RECT 72.870 0.010 72.950 4.280 ;
        RECT 73.790 0.010 73.870 4.280 ;
        RECT 74.710 0.010 74.790 4.280 ;
        RECT 75.630 0.010 75.710 4.280 ;
        RECT 76.550 0.010 76.630 4.280 ;
        RECT 77.470 0.010 77.550 4.280 ;
        RECT 78.390 0.010 78.470 4.280 ;
        RECT 79.310 0.010 79.390 4.280 ;
        RECT 80.230 0.010 80.310 4.280 ;
        RECT 81.150 0.010 81.230 4.280 ;
        RECT 82.070 0.010 82.150 4.280 ;
        RECT 82.990 0.010 83.070 4.280 ;
        RECT 83.910 0.010 83.990 4.280 ;
        RECT 84.830 0.010 84.910 4.280 ;
        RECT 85.750 0.010 85.830 4.280 ;
        RECT 86.670 0.010 86.750 4.280 ;
        RECT 87.590 0.010 87.670 4.280 ;
        RECT 88.510 0.010 88.590 4.280 ;
        RECT 89.430 0.010 89.510 4.280 ;
        RECT 90.350 0.010 90.430 4.280 ;
        RECT 91.270 0.010 91.350 4.280 ;
        RECT 92.190 0.010 92.270 4.280 ;
        RECT 93.110 0.010 93.190 4.280 ;
        RECT 94.030 0.010 94.110 4.280 ;
        RECT 94.950 0.010 95.030 4.280 ;
        RECT 95.870 0.010 95.950 4.280 ;
        RECT 96.790 0.010 199.910 4.280 ;
        RECT 200.750 0.010 200.830 4.280 ;
        RECT 201.670 0.010 201.750 4.280 ;
        RECT 202.590 0.010 202.670 4.280 ;
        RECT 203.510 0.010 203.590 4.280 ;
        RECT 204.430 0.010 204.510 4.280 ;
        RECT 205.350 0.010 205.430 4.280 ;
        RECT 206.270 0.010 206.350 4.280 ;
        RECT 207.190 0.010 207.270 4.280 ;
        RECT 208.110 0.010 208.190 4.280 ;
        RECT 209.030 0.010 209.110 4.280 ;
        RECT 209.950 0.010 210.030 4.280 ;
        RECT 210.870 0.010 210.950 4.280 ;
        RECT 211.790 0.010 211.870 4.280 ;
        RECT 212.710 0.010 212.790 4.280 ;
        RECT 213.630 0.010 213.710 4.280 ;
        RECT 214.550 0.010 214.630 4.280 ;
        RECT 215.470 0.010 215.550 4.280 ;
        RECT 216.390 0.010 216.470 4.280 ;
        RECT 217.310 0.010 217.390 4.280 ;
        RECT 218.230 0.010 218.310 4.280 ;
        RECT 219.150 0.010 219.230 4.280 ;
        RECT 220.070 0.010 220.150 4.280 ;
        RECT 220.990 0.010 221.070 4.280 ;
        RECT 221.910 0.010 221.990 4.280 ;
        RECT 222.830 0.010 222.910 4.280 ;
        RECT 223.750 0.010 223.830 4.280 ;
        RECT 224.670 0.010 224.750 4.280 ;
        RECT 225.590 0.010 225.670 4.280 ;
        RECT 226.510 0.010 226.590 4.280 ;
        RECT 227.430 0.010 227.510 4.280 ;
        RECT 228.350 0.010 228.430 4.280 ;
        RECT 229.270 0.010 229.350 4.280 ;
        RECT 230.190 0.010 230.270 4.280 ;
        RECT 231.110 0.010 231.190 4.280 ;
        RECT 232.030 0.010 232.110 4.280 ;
        RECT 232.950 0.010 233.030 4.280 ;
        RECT 233.870 0.010 233.950 4.280 ;
        RECT 234.790 0.010 234.870 4.280 ;
        RECT 235.710 0.010 235.790 4.280 ;
        RECT 236.630 0.010 236.710 4.280 ;
        RECT 237.550 0.010 237.630 4.280 ;
        RECT 238.470 0.010 238.550 4.280 ;
        RECT 239.390 0.010 239.470 4.280 ;
        RECT 240.310 0.010 240.390 4.280 ;
        RECT 241.230 0.010 241.310 4.280 ;
        RECT 242.150 0.010 242.230 4.280 ;
        RECT 243.070 0.010 243.150 4.280 ;
        RECT 243.990 0.010 244.070 4.280 ;
        RECT 244.910 0.010 244.990 4.280 ;
        RECT 245.830 0.010 245.910 4.280 ;
        RECT 246.750 0.010 246.830 4.280 ;
        RECT 247.670 0.010 247.750 4.280 ;
        RECT 248.590 0.010 248.670 4.280 ;
        RECT 249.510 0.010 249.590 4.280 ;
        RECT 250.430 0.010 250.510 4.280 ;
        RECT 251.350 0.010 251.430 4.280 ;
        RECT 252.270 0.010 252.350 4.280 ;
        RECT 253.190 0.010 253.270 4.280 ;
        RECT 254.110 0.010 254.190 4.280 ;
        RECT 255.030 0.010 255.110 4.280 ;
        RECT 255.950 0.010 256.030 4.280 ;
        RECT 256.870 0.010 256.950 4.280 ;
        RECT 257.790 0.010 257.870 4.280 ;
        RECT 258.710 0.010 258.790 4.280 ;
        RECT 259.630 0.010 259.710 4.280 ;
        RECT 260.550 0.010 260.630 4.280 ;
        RECT 261.470 0.010 261.550 4.280 ;
        RECT 262.390 0.010 262.470 4.280 ;
        RECT 263.310 0.010 263.390 4.280 ;
        RECT 264.230 0.010 264.310 4.280 ;
        RECT 265.150 0.010 265.230 4.280 ;
        RECT 266.070 0.010 266.150 4.280 ;
        RECT 266.990 0.010 267.070 4.280 ;
        RECT 267.910 0.010 267.990 4.280 ;
        RECT 268.830 0.010 268.910 4.280 ;
        RECT 269.750 0.010 269.830 4.280 ;
        RECT 270.670 0.010 270.750 4.280 ;
        RECT 271.590 0.010 271.670 4.280 ;
        RECT 272.510 0.010 272.590 4.280 ;
        RECT 273.430 0.010 273.510 4.280 ;
        RECT 274.350 0.010 274.430 4.280 ;
        RECT 275.270 0.010 275.350 4.280 ;
        RECT 276.190 0.010 276.270 4.280 ;
        RECT 277.110 0.010 277.190 4.280 ;
        RECT 278.030 0.010 278.110 4.280 ;
        RECT 278.950 0.010 279.030 4.280 ;
        RECT 279.870 0.010 279.950 4.280 ;
        RECT 280.790 0.010 280.870 4.280 ;
        RECT 281.710 0.010 281.790 4.280 ;
        RECT 282.630 0.010 282.710 4.280 ;
        RECT 283.550 0.010 283.630 4.280 ;
        RECT 284.470 0.010 284.550 4.280 ;
        RECT 285.390 0.010 285.470 4.280 ;
        RECT 286.310 0.010 286.390 4.280 ;
        RECT 287.230 0.010 287.310 4.280 ;
        RECT 288.150 0.010 288.230 4.280 ;
        RECT 289.070 0.010 289.150 4.280 ;
        RECT 289.990 0.010 290.070 4.280 ;
        RECT 290.910 0.010 290.990 4.280 ;
        RECT 291.830 0.010 291.910 4.280 ;
        RECT 292.750 0.010 292.830 4.280 ;
        RECT 293.670 0.010 293.750 4.280 ;
        RECT 294.590 0.010 294.670 4.280 ;
        RECT 295.510 0.010 295.590 4.280 ;
        RECT 296.430 0.010 699.930 4.280 ;
        RECT 700.770 0.010 700.850 4.280 ;
        RECT 701.690 0.010 701.770 4.280 ;
        RECT 702.610 0.010 702.690 4.280 ;
        RECT 703.530 0.010 703.610 4.280 ;
        RECT 704.450 0.010 704.530 4.280 ;
        RECT 705.370 0.010 705.450 4.280 ;
        RECT 706.290 0.010 706.370 4.280 ;
        RECT 707.210 0.010 707.290 4.280 ;
        RECT 708.130 0.010 708.210 4.280 ;
        RECT 709.050 0.010 709.130 4.280 ;
        RECT 709.970 0.010 710.050 4.280 ;
        RECT 710.890 0.010 710.970 4.280 ;
        RECT 711.810 0.010 711.890 4.280 ;
        RECT 712.730 0.010 712.810 4.280 ;
        RECT 713.650 0.010 713.730 4.280 ;
        RECT 714.570 0.010 714.650 4.280 ;
        RECT 715.490 0.010 715.570 4.280 ;
        RECT 716.410 0.010 716.490 4.280 ;
        RECT 717.330 0.010 717.410 4.280 ;
        RECT 718.250 0.010 718.330 4.280 ;
        RECT 719.170 0.010 719.250 4.280 ;
        RECT 720.090 0.010 720.170 4.280 ;
        RECT 721.010 0.010 721.090 4.280 ;
        RECT 721.930 0.010 722.010 4.280 ;
        RECT 722.850 0.010 722.930 4.280 ;
        RECT 723.770 0.010 723.850 4.280 ;
        RECT 724.690 0.010 724.770 4.280 ;
        RECT 725.610 0.010 725.690 4.280 ;
        RECT 726.530 0.010 726.610 4.280 ;
        RECT 727.450 0.010 727.530 4.280 ;
        RECT 728.370 0.010 728.450 4.280 ;
        RECT 729.290 0.010 729.370 4.280 ;
        RECT 730.210 0.010 730.290 4.280 ;
        RECT 731.130 0.010 731.210 4.280 ;
        RECT 732.050 0.010 732.130 4.280 ;
        RECT 732.970 0.010 733.050 4.280 ;
        RECT 733.890 0.010 733.970 4.280 ;
        RECT 734.810 0.010 734.890 4.280 ;
        RECT 735.730 0.010 735.810 4.280 ;
        RECT 736.650 0.010 736.730 4.280 ;
        RECT 737.570 0.010 737.650 4.280 ;
        RECT 738.490 0.010 738.570 4.280 ;
        RECT 739.410 0.010 739.490 4.280 ;
        RECT 740.330 0.010 740.410 4.280 ;
        RECT 741.250 0.010 741.330 4.280 ;
        RECT 742.170 0.010 742.250 4.280 ;
        RECT 743.090 0.010 743.170 4.280 ;
        RECT 744.010 0.010 744.090 4.280 ;
        RECT 744.930 0.010 745.010 4.280 ;
        RECT 745.850 0.010 745.930 4.280 ;
        RECT 746.770 0.010 746.850 4.280 ;
        RECT 747.690 0.010 747.770 4.280 ;
        RECT 748.610 0.010 748.690 4.280 ;
        RECT 749.530 0.010 749.610 4.280 ;
        RECT 750.450 0.010 750.530 4.280 ;
        RECT 751.370 0.010 751.450 4.280 ;
        RECT 752.290 0.010 752.370 4.280 ;
        RECT 753.210 0.010 753.290 4.280 ;
        RECT 754.130 0.010 754.210 4.280 ;
        RECT 755.050 0.010 755.130 4.280 ;
        RECT 755.970 0.010 756.050 4.280 ;
        RECT 756.890 0.010 756.970 4.280 ;
        RECT 757.810 0.010 757.890 4.280 ;
        RECT 758.730 0.010 758.810 4.280 ;
        RECT 759.650 0.010 759.730 4.280 ;
        RECT 760.570 0.010 760.650 4.280 ;
        RECT 761.490 0.010 761.570 4.280 ;
        RECT 762.410 0.010 762.490 4.280 ;
        RECT 763.330 0.010 763.410 4.280 ;
        RECT 764.250 0.010 764.330 4.280 ;
        RECT 765.170 0.010 765.250 4.280 ;
        RECT 766.090 0.010 766.170 4.280 ;
        RECT 767.010 0.010 767.090 4.280 ;
        RECT 767.930 0.010 768.010 4.280 ;
        RECT 768.850 0.010 768.930 4.280 ;
        RECT 769.770 0.010 769.850 4.280 ;
        RECT 770.690 0.010 770.770 4.280 ;
        RECT 771.610 0.010 771.690 4.280 ;
        RECT 772.530 0.010 772.610 4.280 ;
        RECT 773.450 0.010 773.530 4.280 ;
        RECT 774.370 0.010 774.450 4.280 ;
        RECT 775.290 0.010 775.370 4.280 ;
        RECT 776.210 0.010 776.290 4.280 ;
        RECT 777.130 0.010 777.210 4.280 ;
        RECT 778.050 0.010 778.130 4.280 ;
        RECT 778.970 0.010 779.050 4.280 ;
        RECT 779.890 0.010 779.970 4.280 ;
        RECT 780.810 0.010 780.890 4.280 ;
        RECT 781.730 0.010 781.810 4.280 ;
        RECT 782.650 0.010 782.730 4.280 ;
        RECT 783.570 0.010 783.650 4.280 ;
        RECT 784.490 0.010 784.570 4.280 ;
        RECT 785.410 0.010 785.490 4.280 ;
        RECT 786.330 0.010 786.410 4.280 ;
        RECT 787.250 0.010 787.330 4.280 ;
        RECT 788.170 0.010 788.250 4.280 ;
        RECT 789.090 0.010 789.170 4.280 ;
        RECT 790.010 0.010 790.090 4.280 ;
        RECT 790.930 0.010 791.010 4.280 ;
        RECT 791.850 0.010 791.930 4.280 ;
        RECT 792.770 0.010 792.850 4.280 ;
        RECT 793.690 0.010 793.770 4.280 ;
        RECT 794.610 0.010 794.690 4.280 ;
        RECT 795.530 0.010 795.610 4.280 ;
        RECT 796.450 0.010 1900.070 4.280 ;
        RECT 1900.910 0.010 1900.990 4.280 ;
        RECT 1901.830 0.010 1901.910 4.280 ;
        RECT 1902.750 0.010 1902.830 4.280 ;
        RECT 1903.670 0.010 1903.750 4.280 ;
        RECT 1904.590 0.010 1904.670 4.280 ;
        RECT 1905.510 0.010 1905.590 4.280 ;
        RECT 1906.430 0.010 1906.510 4.280 ;
        RECT 1907.350 0.010 1907.430 4.280 ;
        RECT 1908.270 0.010 1908.350 4.280 ;
        RECT 1909.190 0.010 1909.270 4.280 ;
        RECT 1910.110 0.010 1910.190 4.280 ;
        RECT 1911.030 0.010 1911.110 4.280 ;
        RECT 1911.950 0.010 1912.030 4.280 ;
        RECT 1912.870 0.010 1912.950 4.280 ;
        RECT 1913.790 0.010 1913.870 4.280 ;
        RECT 1914.710 0.010 1914.790 4.280 ;
        RECT 1915.630 0.010 1915.710 4.280 ;
        RECT 1916.550 0.010 1916.630 4.280 ;
        RECT 1917.470 0.010 1917.550 4.280 ;
        RECT 1918.390 0.010 1918.470 4.280 ;
        RECT 1919.310 0.010 1919.390 4.280 ;
        RECT 1920.230 0.010 1920.310 4.280 ;
        RECT 1921.150 0.010 1921.230 4.280 ;
        RECT 1922.070 0.010 1922.150 4.280 ;
        RECT 1922.990 0.010 1923.070 4.280 ;
        RECT 1923.910 0.010 1923.990 4.280 ;
        RECT 1924.830 0.010 1924.910 4.280 ;
        RECT 1925.750 0.010 1925.830 4.280 ;
        RECT 1926.670 0.010 1926.750 4.280 ;
        RECT 1927.590 0.010 1927.670 4.280 ;
        RECT 1928.510 0.010 1928.590 4.280 ;
        RECT 1929.430 0.010 1929.510 4.280 ;
        RECT 1930.350 0.010 1930.430 4.280 ;
        RECT 1931.270 0.010 1931.350 4.280 ;
        RECT 1932.190 0.010 1932.270 4.280 ;
        RECT 1933.110 0.010 1933.190 4.280 ;
        RECT 1934.030 0.010 1934.110 4.280 ;
        RECT 1934.950 0.010 1935.030 4.280 ;
        RECT 1935.870 0.010 1935.950 4.280 ;
        RECT 1936.790 0.010 1936.870 4.280 ;
        RECT 1937.710 0.010 1937.790 4.280 ;
        RECT 1938.630 0.010 1938.710 4.280 ;
        RECT 1939.550 0.010 1939.630 4.280 ;
        RECT 1940.470 0.010 1940.550 4.280 ;
        RECT 1941.390 0.010 1941.470 4.280 ;
        RECT 1942.310 0.010 1942.390 4.280 ;
        RECT 1943.230 0.010 1943.310 4.280 ;
        RECT 1944.150 0.010 1944.230 4.280 ;
        RECT 1945.070 0.010 1945.150 4.280 ;
        RECT 1945.990 0.010 1946.070 4.280 ;
        RECT 1946.910 0.010 1946.990 4.280 ;
        RECT 1947.830 0.010 1947.910 4.280 ;
        RECT 1948.750 0.010 1948.830 4.280 ;
        RECT 1949.670 0.010 1949.750 4.280 ;
        RECT 1950.590 0.010 1950.670 4.280 ;
        RECT 1951.510 0.010 1951.590 4.280 ;
        RECT 1952.430 0.010 1952.510 4.280 ;
        RECT 1953.350 0.010 1953.430 4.280 ;
        RECT 1954.270 0.010 1954.350 4.280 ;
        RECT 1955.190 0.010 1955.270 4.280 ;
        RECT 1956.110 0.010 1956.190 4.280 ;
        RECT 1957.030 0.010 1957.110 4.280 ;
        RECT 1957.950 0.010 1958.030 4.280 ;
        RECT 1958.870 0.010 1958.950 4.280 ;
        RECT 1959.790 0.010 1959.870 4.280 ;
        RECT 1960.710 0.010 1960.790 4.280 ;
        RECT 1961.630 0.010 1961.710 4.280 ;
        RECT 1962.550 0.010 1962.630 4.280 ;
        RECT 1963.470 0.010 1963.550 4.280 ;
        RECT 1964.390 0.010 1964.470 4.280 ;
        RECT 1965.310 0.010 1965.390 4.280 ;
        RECT 1966.230 0.010 1966.310 4.280 ;
        RECT 1967.150 0.010 1967.230 4.280 ;
        RECT 1968.070 0.010 1968.150 4.280 ;
        RECT 1968.990 0.010 1969.070 4.280 ;
        RECT 1969.910 0.010 1969.990 4.280 ;
        RECT 1970.830 0.010 1970.910 4.280 ;
        RECT 1971.750 0.010 1971.830 4.280 ;
        RECT 1972.670 0.010 1972.750 4.280 ;
        RECT 1973.590 0.010 2178.010 4.280 ;
      LAYER met3 ;
        RECT 0.525 3.080 2196.000 145.345 ;
        RECT 0.525 0.320 2195.600 3.080 ;
        RECT 0.525 0.175 2196.000 0.320 ;
      LAYER met4 ;
        RECT 737.075 10.640 1098.100 138.960 ;
        RECT 1101.900 10.640 1462.925 138.960 ;
        RECT 1466.725 10.640 1827.755 138.960 ;
  END
END wb_interconnect
MACRO uart_i2c_usb_spi_top
  CLASS BLOCK ;
  FOREIGN uart_i2c_usb_spi_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 700.000 ;
  PIN app_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 -4.000 0.830 4.000 ;
    END
  END app_clk
  PIN i2c_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 -4.000 73.510 4.000 ;
    END
  END i2c_rstn
  PIN i2cm_intr_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 -4.000 87.310 4.000 ;
    END
  END i2cm_intr_o
  PIN reg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 -4.000 71.670 4.000 ;
    END
  END reg_ack
  PIN reg_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 -4.000 10.950 4.000 ;
    END
  END reg_addr[0]
  PIN reg_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 -4.000 10.030 4.000 ;
    END
  END reg_addr[1]
  PIN reg_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 -4.000 9.110 4.000 ;
    END
  END reg_addr[2]
  PIN reg_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 -4.000 8.190 4.000 ;
    END
  END reg_addr[3]
  PIN reg_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 -4.000 7.270 4.000 ;
    END
  END reg_addr[4]
  PIN reg_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 -4.000 6.350 4.000 ;
    END
  END reg_addr[5]
  PIN reg_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 -4.000 5.430 4.000 ;
    END
  END reg_addr[6]
  PIN reg_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 -4.000 4.510 4.000 ;
    END
  END reg_addr[7]
  PIN reg_be
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 -4.000 11.870 4.000 ;
    END
  END reg_be
  PIN reg_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 -4.000 2.670 4.000 ;
    END
  END reg_cs
  PIN reg_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 -4.000 70.750 4.000 ;
    END
  END reg_rdata[0]
  PIN reg_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 -4.000 61.550 4.000 ;
    END
  END reg_rdata[10]
  PIN reg_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 -4.000 60.630 4.000 ;
    END
  END reg_rdata[11]
  PIN reg_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 -4.000 59.710 4.000 ;
    END
  END reg_rdata[12]
  PIN reg_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 -4.000 58.790 4.000 ;
    END
  END reg_rdata[13]
  PIN reg_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 -4.000 57.870 4.000 ;
    END
  END reg_rdata[14]
  PIN reg_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 -4.000 56.950 4.000 ;
    END
  END reg_rdata[15]
  PIN reg_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 -4.000 56.030 4.000 ;
    END
  END reg_rdata[16]
  PIN reg_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 -4.000 55.110 4.000 ;
    END
  END reg_rdata[17]
  PIN reg_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 -4.000 54.190 4.000 ;
    END
  END reg_rdata[18]
  PIN reg_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 -4.000 53.270 4.000 ;
    END
  END reg_rdata[19]
  PIN reg_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 -4.000 69.830 4.000 ;
    END
  END reg_rdata[1]
  PIN reg_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 -4.000 52.350 4.000 ;
    END
  END reg_rdata[20]
  PIN reg_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 -4.000 51.430 4.000 ;
    END
  END reg_rdata[21]
  PIN reg_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 -4.000 50.510 4.000 ;
    END
  END reg_rdata[22]
  PIN reg_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 -4.000 49.590 4.000 ;
    END
  END reg_rdata[23]
  PIN reg_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 -4.000 48.670 4.000 ;
    END
  END reg_rdata[24]
  PIN reg_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 -4.000 47.750 4.000 ;
    END
  END reg_rdata[25]
  PIN reg_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 -4.000 46.830 4.000 ;
    END
  END reg_rdata[26]
  PIN reg_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 -4.000 45.910 4.000 ;
    END
  END reg_rdata[27]
  PIN reg_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 -4.000 44.990 4.000 ;
    END
  END reg_rdata[28]
  PIN reg_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 -4.000 44.070 4.000 ;
    END
  END reg_rdata[29]
  PIN reg_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 -4.000 68.910 4.000 ;
    END
  END reg_rdata[2]
  PIN reg_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 -4.000 43.150 4.000 ;
    END
  END reg_rdata[30]
  PIN reg_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 -4.000 42.230 4.000 ;
    END
  END reg_rdata[31]
  PIN reg_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 -4.000 67.990 4.000 ;
    END
  END reg_rdata[3]
  PIN reg_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 -4.000 67.070 4.000 ;
    END
  END reg_rdata[4]
  PIN reg_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 -4.000 66.150 4.000 ;
    END
  END reg_rdata[5]
  PIN reg_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 -4.000 65.230 4.000 ;
    END
  END reg_rdata[6]
  PIN reg_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 -4.000 64.310 4.000 ;
    END
  END reg_rdata[7]
  PIN reg_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 -4.000 63.390 4.000 ;
    END
  END reg_rdata[8]
  PIN reg_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 -4.000 62.470 4.000 ;
    END
  END reg_rdata[9]
  PIN reg_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 -4.000 41.310 4.000 ;
    END
  END reg_wdata[0]
  PIN reg_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 -4.000 32.110 4.000 ;
    END
  END reg_wdata[10]
  PIN reg_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 -4.000 31.190 4.000 ;
    END
  END reg_wdata[11]
  PIN reg_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 -4.000 30.270 4.000 ;
    END
  END reg_wdata[12]
  PIN reg_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 -4.000 29.350 4.000 ;
    END
  END reg_wdata[13]
  PIN reg_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 -4.000 28.430 4.000 ;
    END
  END reg_wdata[14]
  PIN reg_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 -4.000 27.510 4.000 ;
    END
  END reg_wdata[15]
  PIN reg_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 -4.000 26.590 4.000 ;
    END
  END reg_wdata[16]
  PIN reg_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 -4.000 25.670 4.000 ;
    END
  END reg_wdata[17]
  PIN reg_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 -4.000 24.750 4.000 ;
    END
  END reg_wdata[18]
  PIN reg_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 -4.000 23.830 4.000 ;
    END
  END reg_wdata[19]
  PIN reg_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 -4.000 40.390 4.000 ;
    END
  END reg_wdata[1]
  PIN reg_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 -4.000 22.910 4.000 ;
    END
  END reg_wdata[20]
  PIN reg_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 -4.000 21.990 4.000 ;
    END
  END reg_wdata[21]
  PIN reg_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 -4.000 21.070 4.000 ;
    END
  END reg_wdata[22]
  PIN reg_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 -4.000 20.150 4.000 ;
    END
  END reg_wdata[23]
  PIN reg_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 -4.000 19.230 4.000 ;
    END
  END reg_wdata[24]
  PIN reg_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 -4.000 18.310 4.000 ;
    END
  END reg_wdata[25]
  PIN reg_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 -4.000 17.390 4.000 ;
    END
  END reg_wdata[26]
  PIN reg_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 -4.000 16.470 4.000 ;
    END
  END reg_wdata[27]
  PIN reg_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 -4.000 15.550 4.000 ;
    END
  END reg_wdata[28]
  PIN reg_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 -4.000 14.630 4.000 ;
    END
  END reg_wdata[29]
  PIN reg_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 -4.000 39.470 4.000 ;
    END
  END reg_wdata[2]
  PIN reg_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 -4.000 13.710 4.000 ;
    END
  END reg_wdata[30]
  PIN reg_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 -4.000 12.790 4.000 ;
    END
  END reg_wdata[31]
  PIN reg_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 -4.000 38.550 4.000 ;
    END
  END reg_wdata[3]
  PIN reg_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 -4.000 37.630 4.000 ;
    END
  END reg_wdata[4]
  PIN reg_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 -4.000 36.710 4.000 ;
    END
  END reg_wdata[5]
  PIN reg_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 -4.000 35.790 4.000 ;
    END
  END reg_wdata[6]
  PIN reg_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 -4.000 34.870 4.000 ;
    END
  END reg_wdata[7]
  PIN reg_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 -4.000 33.950 4.000 ;
    END
  END reg_wdata[8]
  PIN reg_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 -4.000 33.030 4.000 ;
    END
  END reg_wdata[9]
  PIN reg_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 -4.000 3.590 4.000 ;
    END
  END reg_wr
  PIN scl_pad_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 -4.000 75.350 4.000 ;
    END
  END scl_pad_i
  PIN scl_pad_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 -4.000 76.270 4.000 ;
    END
  END scl_pad_o
  PIN scl_pad_oen_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 -4.000 77.190 4.000 ;
    END
  END scl_pad_oen_o
  PIN sda_pad_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 -4.000 78.110 4.000 ;
    END
  END sda_pad_i
  PIN sda_pad_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 -4.000 79.030 4.000 ;
    END
  END sda_pad_o
  PIN sda_padoen_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 -4.000 79.950 4.000 ;
    END
  END sda_padoen_o
  PIN spi_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 -4.000 89.150 4.000 ;
    END
  END spi_rstn
  PIN sspim_sck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 -4.000 90.070 4.000 ;
    END
  END sspim_sck
  PIN sspim_si
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 -4.000 90.990 4.000 ;
    END
  END sspim_si
  PIN sspim_so
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 -4.000 91.910 4.000 ;
    END
  END sspim_so
  PIN sspim_ssn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 -4.000 92.830 4.000 ;
    END
  END sspim_ssn
  PIN uart_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 -4.000 72.590 4.000 ;
    END
  END uart_rstn
  PIN uart_rxd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 -4.000 80.870 4.000 ;
    END
  END uart_rxd
  PIN uart_txd
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 -4.000 81.790 4.000 ;
    END
  END uart_txd
  PIN usb_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 -4.000 1.750 4.000 ;
    END
  END usb_clk
  PIN usb_in_dn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 -4.000 83.630 4.000 ;
    END
  END usb_in_dn
  PIN usb_in_dp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 -4.000 82.710 4.000 ;
    END
  END usb_in_dp
  PIN usb_intr_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 -4.000 88.230 4.000 ;
    END
  END usb_intr_o
  PIN usb_out_dn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 -4.000 85.470 4.000 ;
    END
  END usb_out_dn
  PIN usb_out_dp
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 -4.000 84.550 4.000 ;
    END
  END usb_out_dp
  PIN usb_out_tx_oen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 -4.000 86.390 4.000 ;
    END
  END usb_out_tx_oen
  PIN usb_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 -4.000 74.430 4.000 ;
    END
  END usb_rstn
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.340 10.640 24.340 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.340 10.640 124.340 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 219.340 10.640 224.340 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 319.340 10.640 324.340 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 419.340 10.640 424.340 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 519.340 10.640 524.340 688.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 69.340 10.640 74.340 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 169.340 10.640 174.340 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 269.340 10.640 274.340 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 369.340 10.640 374.340 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 469.340 10.640 474.340 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 569.340 10.640 574.340 688.400 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 4.285 4.845 594.320 688.245 ;
      LAYER met1 ;
        RECT 0.070 0.040 594.320 688.400 ;
      LAYER met2 ;
        RECT 0.100 4.280 591.000 688.400 ;
        RECT 0.100 0.010 0.270 4.280 ;
        RECT 1.110 0.010 1.190 4.280 ;
        RECT 2.030 0.010 2.110 4.280 ;
        RECT 2.950 0.010 3.030 4.280 ;
        RECT 3.870 0.010 3.950 4.280 ;
        RECT 4.790 0.010 4.870 4.280 ;
        RECT 5.710 0.010 5.790 4.280 ;
        RECT 6.630 0.010 6.710 4.280 ;
        RECT 7.550 0.010 7.630 4.280 ;
        RECT 8.470 0.010 8.550 4.280 ;
        RECT 9.390 0.010 9.470 4.280 ;
        RECT 10.310 0.010 10.390 4.280 ;
        RECT 11.230 0.010 11.310 4.280 ;
        RECT 12.150 0.010 12.230 4.280 ;
        RECT 13.070 0.010 13.150 4.280 ;
        RECT 13.990 0.010 14.070 4.280 ;
        RECT 14.910 0.010 14.990 4.280 ;
        RECT 15.830 0.010 15.910 4.280 ;
        RECT 16.750 0.010 16.830 4.280 ;
        RECT 17.670 0.010 17.750 4.280 ;
        RECT 18.590 0.010 18.670 4.280 ;
        RECT 19.510 0.010 19.590 4.280 ;
        RECT 20.430 0.010 20.510 4.280 ;
        RECT 21.350 0.010 21.430 4.280 ;
        RECT 22.270 0.010 22.350 4.280 ;
        RECT 23.190 0.010 23.270 4.280 ;
        RECT 24.110 0.010 24.190 4.280 ;
        RECT 25.030 0.010 25.110 4.280 ;
        RECT 25.950 0.010 26.030 4.280 ;
        RECT 26.870 0.010 26.950 4.280 ;
        RECT 27.790 0.010 27.870 4.280 ;
        RECT 28.710 0.010 28.790 4.280 ;
        RECT 29.630 0.010 29.710 4.280 ;
        RECT 30.550 0.010 30.630 4.280 ;
        RECT 31.470 0.010 31.550 4.280 ;
        RECT 32.390 0.010 32.470 4.280 ;
        RECT 33.310 0.010 33.390 4.280 ;
        RECT 34.230 0.010 34.310 4.280 ;
        RECT 35.150 0.010 35.230 4.280 ;
        RECT 36.070 0.010 36.150 4.280 ;
        RECT 36.990 0.010 37.070 4.280 ;
        RECT 37.910 0.010 37.990 4.280 ;
        RECT 38.830 0.010 38.910 4.280 ;
        RECT 39.750 0.010 39.830 4.280 ;
        RECT 40.670 0.010 40.750 4.280 ;
        RECT 41.590 0.010 41.670 4.280 ;
        RECT 42.510 0.010 42.590 4.280 ;
        RECT 43.430 0.010 43.510 4.280 ;
        RECT 44.350 0.010 44.430 4.280 ;
        RECT 45.270 0.010 45.350 4.280 ;
        RECT 46.190 0.010 46.270 4.280 ;
        RECT 47.110 0.010 47.190 4.280 ;
        RECT 48.030 0.010 48.110 4.280 ;
        RECT 48.950 0.010 49.030 4.280 ;
        RECT 49.870 0.010 49.950 4.280 ;
        RECT 50.790 0.010 50.870 4.280 ;
        RECT 51.710 0.010 51.790 4.280 ;
        RECT 52.630 0.010 52.710 4.280 ;
        RECT 53.550 0.010 53.630 4.280 ;
        RECT 54.470 0.010 54.550 4.280 ;
        RECT 55.390 0.010 55.470 4.280 ;
        RECT 56.310 0.010 56.390 4.280 ;
        RECT 57.230 0.010 57.310 4.280 ;
        RECT 58.150 0.010 58.230 4.280 ;
        RECT 59.070 0.010 59.150 4.280 ;
        RECT 59.990 0.010 60.070 4.280 ;
        RECT 60.910 0.010 60.990 4.280 ;
        RECT 61.830 0.010 61.910 4.280 ;
        RECT 62.750 0.010 62.830 4.280 ;
        RECT 63.670 0.010 63.750 4.280 ;
        RECT 64.590 0.010 64.670 4.280 ;
        RECT 65.510 0.010 65.590 4.280 ;
        RECT 66.430 0.010 66.510 4.280 ;
        RECT 67.350 0.010 67.430 4.280 ;
        RECT 68.270 0.010 68.350 4.280 ;
        RECT 69.190 0.010 69.270 4.280 ;
        RECT 70.110 0.010 70.190 4.280 ;
        RECT 71.030 0.010 71.110 4.280 ;
        RECT 71.950 0.010 72.030 4.280 ;
        RECT 72.870 0.010 72.950 4.280 ;
        RECT 73.790 0.010 73.870 4.280 ;
        RECT 74.710 0.010 74.790 4.280 ;
        RECT 75.630 0.010 75.710 4.280 ;
        RECT 76.550 0.010 76.630 4.280 ;
        RECT 77.470 0.010 77.550 4.280 ;
        RECT 78.390 0.010 78.470 4.280 ;
        RECT 79.310 0.010 79.390 4.280 ;
        RECT 80.230 0.010 80.310 4.280 ;
        RECT 81.150 0.010 81.230 4.280 ;
        RECT 82.070 0.010 82.150 4.280 ;
        RECT 82.990 0.010 83.070 4.280 ;
        RECT 83.910 0.010 83.990 4.280 ;
        RECT 84.830 0.010 84.910 4.280 ;
        RECT 85.750 0.010 85.830 4.280 ;
        RECT 86.670 0.010 86.750 4.280 ;
        RECT 87.590 0.010 87.670 4.280 ;
        RECT 88.510 0.010 88.590 4.280 ;
        RECT 89.430 0.010 89.510 4.280 ;
        RECT 90.350 0.010 90.430 4.280 ;
        RECT 91.270 0.010 91.350 4.280 ;
        RECT 92.190 0.010 92.270 4.280 ;
        RECT 93.110 0.010 591.000 4.280 ;
      LAYER met3 ;
        RECT 1.905 0.175 578.615 688.325 ;
      LAYER met4 ;
        RECT 8.575 10.240 18.940 627.465 ;
        RECT 24.740 10.240 68.940 627.465 ;
        RECT 74.740 10.240 118.940 627.465 ;
        RECT 124.740 10.240 168.940 627.465 ;
        RECT 174.740 10.240 218.940 627.465 ;
        RECT 224.740 10.240 268.940 627.465 ;
        RECT 274.740 10.240 318.940 627.465 ;
        RECT 324.740 10.240 368.940 627.465 ;
        RECT 374.740 10.240 418.940 627.465 ;
        RECT 424.740 10.240 468.940 627.465 ;
        RECT 474.740 10.240 518.585 627.465 ;
        RECT 8.575 1.535 518.585 10.240 ;
  END
END uart_i2c_usb_spi_top
MACRO wb_host
  CLASS BLOCK ;
  FOREIGN wb_host ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 200.000 ;
  PIN cfg_clk_ctrl1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 196.000 114.910 204.000 ;
    END
  END cfg_clk_ctrl1[0]
  PIN cfg_clk_ctrl1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 -4.000 202.310 4.000 ;
    END
  END cfg_clk_ctrl1[10]
  PIN cfg_clk_ctrl1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 -4.000 200.470 4.000 ;
    END
  END cfg_clk_ctrl1[11]
  PIN cfg_clk_ctrl1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 19.760 4.000 20.360 ;
    END
  END cfg_clk_ctrl1[12]
  PIN cfg_clk_ctrl1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 17.040 4.000 17.640 ;
    END
  END cfg_clk_ctrl1[13]
  PIN cfg_clk_ctrl1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 14.320 4.000 14.920 ;
    END
  END cfg_clk_ctrl1[14]
  PIN cfg_clk_ctrl1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 11.600 4.000 12.200 ;
    END
  END cfg_clk_ctrl1[15]
  PIN cfg_clk_ctrl1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 196.000 107.550 204.000 ;
    END
  END cfg_clk_ctrl1[16]
  PIN cfg_clk_ctrl1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 196.000 106.630 204.000 ;
    END
  END cfg_clk_ctrl1[17]
  PIN cfg_clk_ctrl1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 196.000 105.710 204.000 ;
    END
  END cfg_clk_ctrl1[18]
  PIN cfg_clk_ctrl1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 196.000 104.790 204.000 ;
    END
  END cfg_clk_ctrl1[19]
  PIN cfg_clk_ctrl1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 196.000 113.990 204.000 ;
    END
  END cfg_clk_ctrl1[1]
  PIN cfg_clk_ctrl1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 196.000 103.870 204.000 ;
    END
  END cfg_clk_ctrl1[20]
  PIN cfg_clk_ctrl1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 196.000 102.950 204.000 ;
    END
  END cfg_clk_ctrl1[21]
  PIN cfg_clk_ctrl1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 196.000 102.030 204.000 ;
    END
  END cfg_clk_ctrl1[22]
  PIN cfg_clk_ctrl1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 196.000 101.110 204.000 ;
    END
  END cfg_clk_ctrl1[23]
  PIN cfg_clk_ctrl1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 -4.000 213.350 4.000 ;
    END
  END cfg_clk_ctrl1[24]
  PIN cfg_clk_ctrl1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 -4.000 211.510 4.000 ;
    END
  END cfg_clk_ctrl1[25]
  PIN cfg_clk_ctrl1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 -4.000 209.670 4.000 ;
    END
  END cfg_clk_ctrl1[26]
  PIN cfg_clk_ctrl1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 -4.000 207.830 4.000 ;
    END
  END cfg_clk_ctrl1[27]
  PIN cfg_clk_ctrl1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 196.000 100.190 204.000 ;
    END
  END cfg_clk_ctrl1[28]
  PIN cfg_clk_ctrl1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 196.000 99.270 204.000 ;
    END
  END cfg_clk_ctrl1[29]
  PIN cfg_clk_ctrl1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 196.000 113.070 204.000 ;
    END
  END cfg_clk_ctrl1[2]
  PIN cfg_clk_ctrl1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 196.000 98.350 204.000 ;
    END
  END cfg_clk_ctrl1[30]
  PIN cfg_clk_ctrl1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 196.000 97.430 204.000 ;
    END
  END cfg_clk_ctrl1[31]
  PIN cfg_clk_ctrl1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 196.000 112.150 204.000 ;
    END
  END cfg_clk_ctrl1[3]
  PIN cfg_clk_ctrl1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 196.000 111.230 204.000 ;
    END
  END cfg_clk_ctrl1[4]
  PIN cfg_clk_ctrl1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 196.000 110.310 204.000 ;
    END
  END cfg_clk_ctrl1[5]
  PIN cfg_clk_ctrl1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 196.000 109.390 204.000 ;
    END
  END cfg_clk_ctrl1[6]
  PIN cfg_clk_ctrl1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 196.000 108.470 204.000 ;
    END
  END cfg_clk_ctrl1[7]
  PIN cfg_clk_ctrl1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 -4.000 205.990 4.000 ;
    END
  END cfg_clk_ctrl1[8]
  PIN cfg_clk_ctrl1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 -4.000 204.150 4.000 ;
    END
  END cfg_clk_ctrl1[9]
  PIN cfg_clk_ctrl2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 196.000 144.350 204.000 ;
    END
  END cfg_clk_ctrl2[0]
  PIN cfg_clk_ctrl2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 196.000 135.150 204.000 ;
    END
  END cfg_clk_ctrl2[10]
  PIN cfg_clk_ctrl2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 196.000 134.230 204.000 ;
    END
  END cfg_clk_ctrl2[11]
  PIN cfg_clk_ctrl2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 196.000 133.310 204.000 ;
    END
  END cfg_clk_ctrl2[12]
  PIN cfg_clk_ctrl2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 196.000 132.390 204.000 ;
    END
  END cfg_clk_ctrl2[13]
  PIN cfg_clk_ctrl2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 196.000 131.470 204.000 ;
    END
  END cfg_clk_ctrl2[14]
  PIN cfg_clk_ctrl2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 196.000 130.550 204.000 ;
    END
  END cfg_clk_ctrl2[15]
  PIN cfg_clk_ctrl2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 196.000 129.630 204.000 ;
    END
  END cfg_clk_ctrl2[16]
  PIN cfg_clk_ctrl2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 196.000 128.710 204.000 ;
    END
  END cfg_clk_ctrl2[17]
  PIN cfg_clk_ctrl2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 196.000 127.790 204.000 ;
    END
  END cfg_clk_ctrl2[18]
  PIN cfg_clk_ctrl2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 196.000 126.870 204.000 ;
    END
  END cfg_clk_ctrl2[19]
  PIN cfg_clk_ctrl2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 196.000 143.430 204.000 ;
    END
  END cfg_clk_ctrl2[1]
  PIN cfg_clk_ctrl2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 196.000 125.950 204.000 ;
    END
  END cfg_clk_ctrl2[20]
  PIN cfg_clk_ctrl2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 196.000 125.030 204.000 ;
    END
  END cfg_clk_ctrl2[21]
  PIN cfg_clk_ctrl2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 196.000 124.110 204.000 ;
    END
  END cfg_clk_ctrl2[22]
  PIN cfg_clk_ctrl2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 196.000 123.190 204.000 ;
    END
  END cfg_clk_ctrl2[23]
  PIN cfg_clk_ctrl2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 196.000 122.270 204.000 ;
    END
  END cfg_clk_ctrl2[24]
  PIN cfg_clk_ctrl2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 196.000 121.350 204.000 ;
    END
  END cfg_clk_ctrl2[25]
  PIN cfg_clk_ctrl2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 196.000 120.430 204.000 ;
    END
  END cfg_clk_ctrl2[26]
  PIN cfg_clk_ctrl2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 196.000 119.510 204.000 ;
    END
  END cfg_clk_ctrl2[27]
  PIN cfg_clk_ctrl2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 196.000 118.590 204.000 ;
    END
  END cfg_clk_ctrl2[28]
  PIN cfg_clk_ctrl2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 196.000 117.670 204.000 ;
    END
  END cfg_clk_ctrl2[29]
  PIN cfg_clk_ctrl2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 196.000 142.510 204.000 ;
    END
  END cfg_clk_ctrl2[2]
  PIN cfg_clk_ctrl2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 196.000 116.750 204.000 ;
    END
  END cfg_clk_ctrl2[30]
  PIN cfg_clk_ctrl2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 196.000 115.830 204.000 ;
    END
  END cfg_clk_ctrl2[31]
  PIN cfg_clk_ctrl2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 196.000 141.590 204.000 ;
    END
  END cfg_clk_ctrl2[3]
  PIN cfg_clk_ctrl2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 196.000 140.670 204.000 ;
    END
  END cfg_clk_ctrl2[4]
  PIN cfg_clk_ctrl2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 196.000 139.750 204.000 ;
    END
  END cfg_clk_ctrl2[5]
  PIN cfg_clk_ctrl2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 196.000 138.830 204.000 ;
    END
  END cfg_clk_ctrl2[6]
  PIN cfg_clk_ctrl2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 196.000 137.910 204.000 ;
    END
  END cfg_clk_ctrl2[7]
  PIN cfg_clk_ctrl2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 196.000 136.990 204.000 ;
    END
  END cfg_clk_ctrl2[8]
  PIN cfg_clk_ctrl2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 196.000 136.070 204.000 ;
    END
  END cfg_clk_ctrl2[9]
  PIN cpu_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 -4.000 404.250 4.000 ;
    END
  END cpu_clk
  PIN cpu_rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 6.160 4.000 6.760 ;
    END
  END cpu_rst_n
  PIN i2cm_rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 196.000 146.190 204.000 ;
    END
  END i2cm_rst_n
  PIN qspim_rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 8.880 4.000 9.480 ;
    END
  END qspim_rst_n
  PIN rtc_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 -4.000 406.090 4.000 ;
    END
  END rtc_clk
  PIN sdram_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 0.720 4.000 1.320 ;
    END
  END sdram_clk
  PIN sspim_rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 3.440 4.000 4.040 ;
    END
  END sspim_rst_n
  PIN uart_i2c_usb_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 196.000 149.870 204.000 ;
    END
  END uart_i2c_usb_sel[0]
  PIN uart_i2c_usb_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 196.000 148.950 204.000 ;
    END
  END uart_i2c_usb_sel[1]
  PIN uart_rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 196.000 145.270 204.000 ;
    END
  END uart_rst_n
  PIN usb_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 196.000 148.030 204.000 ;
    END
  END usb_clk
  PIN usb_rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 196.000 147.110 204.000 ;
    END
  END usb_rst_n
  PIN user_clock1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 -4.000 1.750 4.000 ;
    END
  END user_clock1
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 -4.000 0.830 4.000 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.340 10.640 24.340 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.340 10.640 124.340 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 219.340 10.640 224.340 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 319.340 10.640 324.340 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 419.340 10.640 424.340 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 69.340 10.640 74.340 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 169.340 10.640 174.340 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 269.340 10.640 274.340 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 369.340 10.640 374.340 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 469.340 10.640 474.340 187.920 ;
    END
  END vssd1
  PIN wbd_int_rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 196.000 150.790 204.000 ;
    END
  END wbd_int_rst_n
  PIN wbm_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 -4.000 4.510 4.000 ;
    END
  END wbm_ack_o
  PIN wbm_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 -4.000 8.190 4.000 ;
    END
  END wbm_adr_i[0]
  PIN wbm_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 -4.000 39.470 4.000 ;
    END
  END wbm_adr_i[10]
  PIN wbm_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 -4.000 42.230 4.000 ;
    END
  END wbm_adr_i[11]
  PIN wbm_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 -4.000 44.990 4.000 ;
    END
  END wbm_adr_i[12]
  PIN wbm_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 -4.000 47.750 4.000 ;
    END
  END wbm_adr_i[13]
  PIN wbm_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 -4.000 50.510 4.000 ;
    END
  END wbm_adr_i[14]
  PIN wbm_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 -4.000 53.270 4.000 ;
    END
  END wbm_adr_i[15]
  PIN wbm_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 -4.000 56.030 4.000 ;
    END
  END wbm_adr_i[16]
  PIN wbm_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 -4.000 58.790 4.000 ;
    END
  END wbm_adr_i[17]
  PIN wbm_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 -4.000 61.550 4.000 ;
    END
  END wbm_adr_i[18]
  PIN wbm_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 -4.000 64.310 4.000 ;
    END
  END wbm_adr_i[19]
  PIN wbm_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 -4.000 11.870 4.000 ;
    END
  END wbm_adr_i[1]
  PIN wbm_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 -4.000 67.070 4.000 ;
    END
  END wbm_adr_i[20]
  PIN wbm_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 -4.000 69.830 4.000 ;
    END
  END wbm_adr_i[21]
  PIN wbm_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 -4.000 72.590 4.000 ;
    END
  END wbm_adr_i[22]
  PIN wbm_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 -4.000 75.350 4.000 ;
    END
  END wbm_adr_i[23]
  PIN wbm_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 -4.000 78.110 4.000 ;
    END
  END wbm_adr_i[24]
  PIN wbm_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 -4.000 80.870 4.000 ;
    END
  END wbm_adr_i[25]
  PIN wbm_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 -4.000 83.630 4.000 ;
    END
  END wbm_adr_i[26]
  PIN wbm_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 -4.000 86.390 4.000 ;
    END
  END wbm_adr_i[27]
  PIN wbm_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 -4.000 89.150 4.000 ;
    END
  END wbm_adr_i[28]
  PIN wbm_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 -4.000 91.910 4.000 ;
    END
  END wbm_adr_i[29]
  PIN wbm_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 -4.000 15.550 4.000 ;
    END
  END wbm_adr_i[2]
  PIN wbm_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 -4.000 94.670 4.000 ;
    END
  END wbm_adr_i[30]
  PIN wbm_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 -4.000 97.430 4.000 ;
    END
  END wbm_adr_i[31]
  PIN wbm_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 -4.000 19.230 4.000 ;
    END
  END wbm_adr_i[3]
  PIN wbm_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 -4.000 22.910 4.000 ;
    END
  END wbm_adr_i[4]
  PIN wbm_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 -4.000 25.670 4.000 ;
    END
  END wbm_adr_i[5]
  PIN wbm_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 -4.000 28.430 4.000 ;
    END
  END wbm_adr_i[6]
  PIN wbm_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 -4.000 31.190 4.000 ;
    END
  END wbm_adr_i[7]
  PIN wbm_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 -4.000 33.950 4.000 ;
    END
  END wbm_adr_i[8]
  PIN wbm_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 -4.000 36.710 4.000 ;
    END
  END wbm_adr_i[9]
  PIN wbm_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 -4.000 2.670 4.000 ;
    END
  END wbm_clk_i
  PIN wbm_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 -4.000 5.430 4.000 ;
    END
  END wbm_cyc_i
  PIN wbm_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 -4.000 9.110 4.000 ;
    END
  END wbm_dat_i[0]
  PIN wbm_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 -4.000 40.390 4.000 ;
    END
  END wbm_dat_i[10]
  PIN wbm_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 -4.000 43.150 4.000 ;
    END
  END wbm_dat_i[11]
  PIN wbm_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 -4.000 45.910 4.000 ;
    END
  END wbm_dat_i[12]
  PIN wbm_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 -4.000 48.670 4.000 ;
    END
  END wbm_dat_i[13]
  PIN wbm_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 -4.000 51.430 4.000 ;
    END
  END wbm_dat_i[14]
  PIN wbm_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 -4.000 54.190 4.000 ;
    END
  END wbm_dat_i[15]
  PIN wbm_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 -4.000 56.950 4.000 ;
    END
  END wbm_dat_i[16]
  PIN wbm_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 -4.000 59.710 4.000 ;
    END
  END wbm_dat_i[17]
  PIN wbm_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 -4.000 62.470 4.000 ;
    END
  END wbm_dat_i[18]
  PIN wbm_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 -4.000 65.230 4.000 ;
    END
  END wbm_dat_i[19]
  PIN wbm_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 -4.000 12.790 4.000 ;
    END
  END wbm_dat_i[1]
  PIN wbm_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 -4.000 67.990 4.000 ;
    END
  END wbm_dat_i[20]
  PIN wbm_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 -4.000 70.750 4.000 ;
    END
  END wbm_dat_i[21]
  PIN wbm_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 -4.000 73.510 4.000 ;
    END
  END wbm_dat_i[22]
  PIN wbm_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 -4.000 76.270 4.000 ;
    END
  END wbm_dat_i[23]
  PIN wbm_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 -4.000 79.030 4.000 ;
    END
  END wbm_dat_i[24]
  PIN wbm_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 -4.000 81.790 4.000 ;
    END
  END wbm_dat_i[25]
  PIN wbm_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 -4.000 84.550 4.000 ;
    END
  END wbm_dat_i[26]
  PIN wbm_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 -4.000 87.310 4.000 ;
    END
  END wbm_dat_i[27]
  PIN wbm_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 -4.000 90.070 4.000 ;
    END
  END wbm_dat_i[28]
  PIN wbm_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 -4.000 92.830 4.000 ;
    END
  END wbm_dat_i[29]
  PIN wbm_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 -4.000 16.470 4.000 ;
    END
  END wbm_dat_i[2]
  PIN wbm_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 -4.000 95.590 4.000 ;
    END
  END wbm_dat_i[30]
  PIN wbm_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 -4.000 98.350 4.000 ;
    END
  END wbm_dat_i[31]
  PIN wbm_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 -4.000 20.150 4.000 ;
    END
  END wbm_dat_i[3]
  PIN wbm_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 -4.000 23.830 4.000 ;
    END
  END wbm_dat_i[4]
  PIN wbm_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 -4.000 26.590 4.000 ;
    END
  END wbm_dat_i[5]
  PIN wbm_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 -4.000 29.350 4.000 ;
    END
  END wbm_dat_i[6]
  PIN wbm_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 -4.000 32.110 4.000 ;
    END
  END wbm_dat_i[7]
  PIN wbm_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 -4.000 34.870 4.000 ;
    END
  END wbm_dat_i[8]
  PIN wbm_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 -4.000 37.630 4.000 ;
    END
  END wbm_dat_i[9]
  PIN wbm_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 -4.000 10.030 4.000 ;
    END
  END wbm_dat_o[0]
  PIN wbm_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 -4.000 41.310 4.000 ;
    END
  END wbm_dat_o[10]
  PIN wbm_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 -4.000 44.070 4.000 ;
    END
  END wbm_dat_o[11]
  PIN wbm_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 -4.000 46.830 4.000 ;
    END
  END wbm_dat_o[12]
  PIN wbm_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 -4.000 49.590 4.000 ;
    END
  END wbm_dat_o[13]
  PIN wbm_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 -4.000 52.350 4.000 ;
    END
  END wbm_dat_o[14]
  PIN wbm_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 -4.000 55.110 4.000 ;
    END
  END wbm_dat_o[15]
  PIN wbm_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 -4.000 57.870 4.000 ;
    END
  END wbm_dat_o[16]
  PIN wbm_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 -4.000 60.630 4.000 ;
    END
  END wbm_dat_o[17]
  PIN wbm_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 -4.000 63.390 4.000 ;
    END
  END wbm_dat_o[18]
  PIN wbm_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 -4.000 66.150 4.000 ;
    END
  END wbm_dat_o[19]
  PIN wbm_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 -4.000 13.710 4.000 ;
    END
  END wbm_dat_o[1]
  PIN wbm_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 -4.000 68.910 4.000 ;
    END
  END wbm_dat_o[20]
  PIN wbm_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 -4.000 71.670 4.000 ;
    END
  END wbm_dat_o[21]
  PIN wbm_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 -4.000 74.430 4.000 ;
    END
  END wbm_dat_o[22]
  PIN wbm_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 -4.000 77.190 4.000 ;
    END
  END wbm_dat_o[23]
  PIN wbm_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 -4.000 79.950 4.000 ;
    END
  END wbm_dat_o[24]
  PIN wbm_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 -4.000 82.710 4.000 ;
    END
  END wbm_dat_o[25]
  PIN wbm_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 -4.000 85.470 4.000 ;
    END
  END wbm_dat_o[26]
  PIN wbm_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 -4.000 88.230 4.000 ;
    END
  END wbm_dat_o[27]
  PIN wbm_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 -4.000 90.990 4.000 ;
    END
  END wbm_dat_o[28]
  PIN wbm_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 -4.000 93.750 4.000 ;
    END
  END wbm_dat_o[29]
  PIN wbm_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 -4.000 17.390 4.000 ;
    END
  END wbm_dat_o[2]
  PIN wbm_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 -4.000 96.510 4.000 ;
    END
  END wbm_dat_o[30]
  PIN wbm_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 -4.000 99.270 4.000 ;
    END
  END wbm_dat_o[31]
  PIN wbm_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 -4.000 21.070 4.000 ;
    END
  END wbm_dat_o[3]
  PIN wbm_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 -4.000 24.750 4.000 ;
    END
  END wbm_dat_o[4]
  PIN wbm_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 -4.000 27.510 4.000 ;
    END
  END wbm_dat_o[5]
  PIN wbm_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 -4.000 30.270 4.000 ;
    END
  END wbm_dat_o[6]
  PIN wbm_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 -4.000 33.030 4.000 ;
    END
  END wbm_dat_o[7]
  PIN wbm_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 -4.000 35.790 4.000 ;
    END
  END wbm_dat_o[8]
  PIN wbm_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 -4.000 38.550 4.000 ;
    END
  END wbm_dat_o[9]
  PIN wbm_err_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 -4.000 100.190 4.000 ;
    END
  END wbm_err_o
  PIN wbm_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 -4.000 3.590 4.000 ;
    END
  END wbm_rst_i
  PIN wbm_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 -4.000 10.950 4.000 ;
    END
  END wbm_sel_i[0]
  PIN wbm_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 -4.000 14.630 4.000 ;
    END
  END wbm_sel_i[1]
  PIN wbm_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 -4.000 18.310 4.000 ;
    END
  END wbm_sel_i[2]
  PIN wbm_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 -4.000 21.990 4.000 ;
    END
  END wbm_sel_i[3]
  PIN wbm_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 -4.000 6.350 4.000 ;
    END
  END wbm_stb_i
  PIN wbm_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 -4.000 7.270 4.000 ;
    END
  END wbm_we_i
  PIN wbs_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 196.000 94.670 204.000 ;
    END
  END wbs_ack_i
  PIN wbs_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 196.000 31.190 204.000 ;
    END
  END wbs_adr_o[0]
  PIN wbs_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 196.000 21.990 204.000 ;
    END
  END wbs_adr_o[10]
  PIN wbs_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 196.000 21.070 204.000 ;
    END
  END wbs_adr_o[11]
  PIN wbs_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 196.000 20.150 204.000 ;
    END
  END wbs_adr_o[12]
  PIN wbs_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 196.000 19.230 204.000 ;
    END
  END wbs_adr_o[13]
  PIN wbs_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 196.000 18.310 204.000 ;
    END
  END wbs_adr_o[14]
  PIN wbs_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 196.000 17.390 204.000 ;
    END
  END wbs_adr_o[15]
  PIN wbs_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 196.000 16.470 204.000 ;
    END
  END wbs_adr_o[16]
  PIN wbs_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 196.000 15.550 204.000 ;
    END
  END wbs_adr_o[17]
  PIN wbs_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 196.000 14.630 204.000 ;
    END
  END wbs_adr_o[18]
  PIN wbs_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 196.000 13.710 204.000 ;
    END
  END wbs_adr_o[19]
  PIN wbs_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 196.000 30.270 204.000 ;
    END
  END wbs_adr_o[1]
  PIN wbs_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 196.000 12.790 204.000 ;
    END
  END wbs_adr_o[20]
  PIN wbs_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 196.000 11.870 204.000 ;
    END
  END wbs_adr_o[21]
  PIN wbs_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 196.000 10.950 204.000 ;
    END
  END wbs_adr_o[22]
  PIN wbs_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 196.000 10.030 204.000 ;
    END
  END wbs_adr_o[23]
  PIN wbs_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 196.000 9.110 204.000 ;
    END
  END wbs_adr_o[24]
  PIN wbs_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 196.000 8.190 204.000 ;
    END
  END wbs_adr_o[25]
  PIN wbs_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 196.000 7.270 204.000 ;
    END
  END wbs_adr_o[26]
  PIN wbs_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 196.000 6.350 204.000 ;
    END
  END wbs_adr_o[27]
  PIN wbs_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 196.000 5.430 204.000 ;
    END
  END wbs_adr_o[28]
  PIN wbs_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 196.000 4.510 204.000 ;
    END
  END wbs_adr_o[29]
  PIN wbs_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 196.000 29.350 204.000 ;
    END
  END wbs_adr_o[2]
  PIN wbs_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 196.000 3.590 204.000 ;
    END
  END wbs_adr_o[30]
  PIN wbs_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 196.000 2.670 204.000 ;
    END
  END wbs_adr_o[31]
  PIN wbs_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 196.000 28.430 204.000 ;
    END
  END wbs_adr_o[3]
  PIN wbs_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 196.000 27.510 204.000 ;
    END
  END wbs_adr_o[4]
  PIN wbs_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 196.000 26.590 204.000 ;
    END
  END wbs_adr_o[5]
  PIN wbs_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 196.000 25.670 204.000 ;
    END
  END wbs_adr_o[6]
  PIN wbs_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 196.000 24.750 204.000 ;
    END
  END wbs_adr_o[7]
  PIN wbs_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 196.000 23.830 204.000 ;
    END
  END wbs_adr_o[8]
  PIN wbs_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 196.000 22.910 204.000 ;
    END
  END wbs_adr_o[9]
  PIN wbs_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 -4.000 400.570 4.000 ;
    END
  END wbs_clk_i
  PIN wbs_clk_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 -4.000 402.410 4.000 ;
    END
  END wbs_clk_out
  PIN wbs_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 196.000 96.510 204.000 ;
    END
  END wbs_cyc_o
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 196.000 93.750 204.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 196.000 84.550 204.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 196.000 83.630 204.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 196.000 82.710 204.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 196.000 81.790 204.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 196.000 80.870 204.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 196.000 79.950 204.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 196.000 79.030 204.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 196.000 78.110 204.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 196.000 77.190 204.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 196.000 76.270 204.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 196.000 92.830 204.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 196.000 75.350 204.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 196.000 74.430 204.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 196.000 73.510 204.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 196.000 72.590 204.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 196.000 71.670 204.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 196.000 70.750 204.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 196.000 69.830 204.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 196.000 68.910 204.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 196.000 67.990 204.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 196.000 67.070 204.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 196.000 91.910 204.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 196.000 66.150 204.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 196.000 65.230 204.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 196.000 90.990 204.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 196.000 90.070 204.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 196.000 89.150 204.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 196.000 88.230 204.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 196.000 87.310 204.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 196.000 86.390 204.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 196.000 85.470 204.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 196.000 64.310 204.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 196.000 55.110 204.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 196.000 54.190 204.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 196.000 53.270 204.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 196.000 52.350 204.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 196.000 51.430 204.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 196.000 50.510 204.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 196.000 49.590 204.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 196.000 48.670 204.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 196.000 47.750 204.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 196.000 46.830 204.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 196.000 63.390 204.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 196.000 45.910 204.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 196.000 44.990 204.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 196.000 44.070 204.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 196.000 43.150 204.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 196.000 42.230 204.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 196.000 41.310 204.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 196.000 40.390 204.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 196.000 39.470 204.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 196.000 38.550 204.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 196.000 37.630 204.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 196.000 62.470 204.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 196.000 36.710 204.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 196.000 35.790 204.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 196.000 61.550 204.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 196.000 60.630 204.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 196.000 59.710 204.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 196.000 58.790 204.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 196.000 57.870 204.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 196.000 56.950 204.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 196.000 56.030 204.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 196.000 95.590 204.000 ;
    END
  END wbs_err_i
  PIN wbs_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 196.000 34.870 204.000 ;
    END
  END wbs_sel_o[0]
  PIN wbs_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 196.000 33.950 204.000 ;
    END
  END wbs_sel_o[1]
  PIN wbs_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 196.000 33.030 204.000 ;
    END
  END wbs_sel_o[2]
  PIN wbs_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 196.000 32.110 204.000 ;
    END
  END wbs_sel_o[3]
  PIN wbs_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 196.000 0.830 204.000 ;
    END
  END wbs_stb_o
  PIN wbs_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 196.000 1.750 204.000 ;
    END
  END wbs_we_o
  OBS
      LAYER li1 ;
        RECT 4.745 1.445 494.040 198.135 ;
      LAYER met1 ;
        RECT 0.070 0.040 494.040 199.200 ;
      LAYER met2 ;
        RECT 0.100 195.720 0.270 199.230 ;
        RECT 1.110 195.720 1.190 199.230 ;
        RECT 2.030 195.720 2.110 199.230 ;
        RECT 2.950 195.720 3.030 199.230 ;
        RECT 3.870 195.720 3.950 199.230 ;
        RECT 4.790 195.720 4.870 199.230 ;
        RECT 5.710 195.720 5.790 199.230 ;
        RECT 6.630 195.720 6.710 199.230 ;
        RECT 7.550 195.720 7.630 199.230 ;
        RECT 8.470 195.720 8.550 199.230 ;
        RECT 9.390 195.720 9.470 199.230 ;
        RECT 10.310 195.720 10.390 199.230 ;
        RECT 11.230 195.720 11.310 199.230 ;
        RECT 12.150 195.720 12.230 199.230 ;
        RECT 13.070 195.720 13.150 199.230 ;
        RECT 13.990 195.720 14.070 199.230 ;
        RECT 14.910 195.720 14.990 199.230 ;
        RECT 15.830 195.720 15.910 199.230 ;
        RECT 16.750 195.720 16.830 199.230 ;
        RECT 17.670 195.720 17.750 199.230 ;
        RECT 18.590 195.720 18.670 199.230 ;
        RECT 19.510 195.720 19.590 199.230 ;
        RECT 20.430 195.720 20.510 199.230 ;
        RECT 21.350 195.720 21.430 199.230 ;
        RECT 22.270 195.720 22.350 199.230 ;
        RECT 23.190 195.720 23.270 199.230 ;
        RECT 24.110 195.720 24.190 199.230 ;
        RECT 25.030 195.720 25.110 199.230 ;
        RECT 25.950 195.720 26.030 199.230 ;
        RECT 26.870 195.720 26.950 199.230 ;
        RECT 27.790 195.720 27.870 199.230 ;
        RECT 28.710 195.720 28.790 199.230 ;
        RECT 29.630 195.720 29.710 199.230 ;
        RECT 30.550 195.720 30.630 199.230 ;
        RECT 31.470 195.720 31.550 199.230 ;
        RECT 32.390 195.720 32.470 199.230 ;
        RECT 33.310 195.720 33.390 199.230 ;
        RECT 34.230 195.720 34.310 199.230 ;
        RECT 35.150 195.720 35.230 199.230 ;
        RECT 36.070 195.720 36.150 199.230 ;
        RECT 36.990 195.720 37.070 199.230 ;
        RECT 37.910 195.720 37.990 199.230 ;
        RECT 38.830 195.720 38.910 199.230 ;
        RECT 39.750 195.720 39.830 199.230 ;
        RECT 40.670 195.720 40.750 199.230 ;
        RECT 41.590 195.720 41.670 199.230 ;
        RECT 42.510 195.720 42.590 199.230 ;
        RECT 43.430 195.720 43.510 199.230 ;
        RECT 44.350 195.720 44.430 199.230 ;
        RECT 45.270 195.720 45.350 199.230 ;
        RECT 46.190 195.720 46.270 199.230 ;
        RECT 47.110 195.720 47.190 199.230 ;
        RECT 48.030 195.720 48.110 199.230 ;
        RECT 48.950 195.720 49.030 199.230 ;
        RECT 49.870 195.720 49.950 199.230 ;
        RECT 50.790 195.720 50.870 199.230 ;
        RECT 51.710 195.720 51.790 199.230 ;
        RECT 52.630 195.720 52.710 199.230 ;
        RECT 53.550 195.720 53.630 199.230 ;
        RECT 54.470 195.720 54.550 199.230 ;
        RECT 55.390 195.720 55.470 199.230 ;
        RECT 56.310 195.720 56.390 199.230 ;
        RECT 57.230 195.720 57.310 199.230 ;
        RECT 58.150 195.720 58.230 199.230 ;
        RECT 59.070 195.720 59.150 199.230 ;
        RECT 59.990 195.720 60.070 199.230 ;
        RECT 60.910 195.720 60.990 199.230 ;
        RECT 61.830 195.720 61.910 199.230 ;
        RECT 62.750 195.720 62.830 199.230 ;
        RECT 63.670 195.720 63.750 199.230 ;
        RECT 64.590 195.720 64.670 199.230 ;
        RECT 65.510 195.720 65.590 199.230 ;
        RECT 66.430 195.720 66.510 199.230 ;
        RECT 67.350 195.720 67.430 199.230 ;
        RECT 68.270 195.720 68.350 199.230 ;
        RECT 69.190 195.720 69.270 199.230 ;
        RECT 70.110 195.720 70.190 199.230 ;
        RECT 71.030 195.720 71.110 199.230 ;
        RECT 71.950 195.720 72.030 199.230 ;
        RECT 72.870 195.720 72.950 199.230 ;
        RECT 73.790 195.720 73.870 199.230 ;
        RECT 74.710 195.720 74.790 199.230 ;
        RECT 75.630 195.720 75.710 199.230 ;
        RECT 76.550 195.720 76.630 199.230 ;
        RECT 77.470 195.720 77.550 199.230 ;
        RECT 78.390 195.720 78.470 199.230 ;
        RECT 79.310 195.720 79.390 199.230 ;
        RECT 80.230 195.720 80.310 199.230 ;
        RECT 81.150 195.720 81.230 199.230 ;
        RECT 82.070 195.720 82.150 199.230 ;
        RECT 82.990 195.720 83.070 199.230 ;
        RECT 83.910 195.720 83.990 199.230 ;
        RECT 84.830 195.720 84.910 199.230 ;
        RECT 85.750 195.720 85.830 199.230 ;
        RECT 86.670 195.720 86.750 199.230 ;
        RECT 87.590 195.720 87.670 199.230 ;
        RECT 88.510 195.720 88.590 199.230 ;
        RECT 89.430 195.720 89.510 199.230 ;
        RECT 90.350 195.720 90.430 199.230 ;
        RECT 91.270 195.720 91.350 199.230 ;
        RECT 92.190 195.720 92.270 199.230 ;
        RECT 93.110 195.720 93.190 199.230 ;
        RECT 94.030 195.720 94.110 199.230 ;
        RECT 94.950 195.720 95.030 199.230 ;
        RECT 95.870 195.720 95.950 199.230 ;
        RECT 96.790 195.720 96.870 199.230 ;
        RECT 97.710 195.720 97.790 199.230 ;
        RECT 98.630 195.720 98.710 199.230 ;
        RECT 99.550 195.720 99.630 199.230 ;
        RECT 100.470 195.720 100.550 199.230 ;
        RECT 101.390 195.720 101.470 199.230 ;
        RECT 102.310 195.720 102.390 199.230 ;
        RECT 103.230 195.720 103.310 199.230 ;
        RECT 104.150 195.720 104.230 199.230 ;
        RECT 105.070 195.720 105.150 199.230 ;
        RECT 105.990 195.720 106.070 199.230 ;
        RECT 106.910 195.720 106.990 199.230 ;
        RECT 107.830 195.720 107.910 199.230 ;
        RECT 108.750 195.720 108.830 199.230 ;
        RECT 109.670 195.720 109.750 199.230 ;
        RECT 110.590 195.720 110.670 199.230 ;
        RECT 111.510 195.720 111.590 199.230 ;
        RECT 112.430 195.720 112.510 199.230 ;
        RECT 113.350 195.720 113.430 199.230 ;
        RECT 114.270 195.720 114.350 199.230 ;
        RECT 115.190 195.720 115.270 199.230 ;
        RECT 116.110 195.720 116.190 199.230 ;
        RECT 117.030 195.720 117.110 199.230 ;
        RECT 117.950 195.720 118.030 199.230 ;
        RECT 118.870 195.720 118.950 199.230 ;
        RECT 119.790 195.720 119.870 199.230 ;
        RECT 120.710 195.720 120.790 199.230 ;
        RECT 121.630 195.720 121.710 199.230 ;
        RECT 122.550 195.720 122.630 199.230 ;
        RECT 123.470 195.720 123.550 199.230 ;
        RECT 124.390 195.720 124.470 199.230 ;
        RECT 125.310 195.720 125.390 199.230 ;
        RECT 126.230 195.720 126.310 199.230 ;
        RECT 127.150 195.720 127.230 199.230 ;
        RECT 128.070 195.720 128.150 199.230 ;
        RECT 128.990 195.720 129.070 199.230 ;
        RECT 129.910 195.720 129.990 199.230 ;
        RECT 130.830 195.720 130.910 199.230 ;
        RECT 131.750 195.720 131.830 199.230 ;
        RECT 132.670 195.720 132.750 199.230 ;
        RECT 133.590 195.720 133.670 199.230 ;
        RECT 134.510 195.720 134.590 199.230 ;
        RECT 135.430 195.720 135.510 199.230 ;
        RECT 136.350 195.720 136.430 199.230 ;
        RECT 137.270 195.720 137.350 199.230 ;
        RECT 138.190 195.720 138.270 199.230 ;
        RECT 139.110 195.720 139.190 199.230 ;
        RECT 140.030 195.720 140.110 199.230 ;
        RECT 140.950 195.720 141.030 199.230 ;
        RECT 141.870 195.720 141.950 199.230 ;
        RECT 142.790 195.720 142.870 199.230 ;
        RECT 143.710 195.720 143.790 199.230 ;
        RECT 144.630 195.720 144.710 199.230 ;
        RECT 145.550 195.720 145.630 199.230 ;
        RECT 146.470 195.720 146.550 199.230 ;
        RECT 147.390 195.720 147.470 199.230 ;
        RECT 148.310 195.720 148.390 199.230 ;
        RECT 149.230 195.720 149.310 199.230 ;
        RECT 150.150 195.720 150.230 199.230 ;
        RECT 151.070 195.720 474.210 199.230 ;
        RECT 0.100 4.280 474.210 195.720 ;
        RECT 0.100 0.010 0.270 4.280 ;
        RECT 1.110 0.010 1.190 4.280 ;
        RECT 2.030 0.010 2.110 4.280 ;
        RECT 2.950 0.010 3.030 4.280 ;
        RECT 3.870 0.010 3.950 4.280 ;
        RECT 4.790 0.010 4.870 4.280 ;
        RECT 5.710 0.010 5.790 4.280 ;
        RECT 6.630 0.010 6.710 4.280 ;
        RECT 7.550 0.010 7.630 4.280 ;
        RECT 8.470 0.010 8.550 4.280 ;
        RECT 9.390 0.010 9.470 4.280 ;
        RECT 10.310 0.010 10.390 4.280 ;
        RECT 11.230 0.010 11.310 4.280 ;
        RECT 12.150 0.010 12.230 4.280 ;
        RECT 13.070 0.010 13.150 4.280 ;
        RECT 13.990 0.010 14.070 4.280 ;
        RECT 14.910 0.010 14.990 4.280 ;
        RECT 15.830 0.010 15.910 4.280 ;
        RECT 16.750 0.010 16.830 4.280 ;
        RECT 17.670 0.010 17.750 4.280 ;
        RECT 18.590 0.010 18.670 4.280 ;
        RECT 19.510 0.010 19.590 4.280 ;
        RECT 20.430 0.010 20.510 4.280 ;
        RECT 21.350 0.010 21.430 4.280 ;
        RECT 22.270 0.010 22.350 4.280 ;
        RECT 23.190 0.010 23.270 4.280 ;
        RECT 24.110 0.010 24.190 4.280 ;
        RECT 25.030 0.010 25.110 4.280 ;
        RECT 25.950 0.010 26.030 4.280 ;
        RECT 26.870 0.010 26.950 4.280 ;
        RECT 27.790 0.010 27.870 4.280 ;
        RECT 28.710 0.010 28.790 4.280 ;
        RECT 29.630 0.010 29.710 4.280 ;
        RECT 30.550 0.010 30.630 4.280 ;
        RECT 31.470 0.010 31.550 4.280 ;
        RECT 32.390 0.010 32.470 4.280 ;
        RECT 33.310 0.010 33.390 4.280 ;
        RECT 34.230 0.010 34.310 4.280 ;
        RECT 35.150 0.010 35.230 4.280 ;
        RECT 36.070 0.010 36.150 4.280 ;
        RECT 36.990 0.010 37.070 4.280 ;
        RECT 37.910 0.010 37.990 4.280 ;
        RECT 38.830 0.010 38.910 4.280 ;
        RECT 39.750 0.010 39.830 4.280 ;
        RECT 40.670 0.010 40.750 4.280 ;
        RECT 41.590 0.010 41.670 4.280 ;
        RECT 42.510 0.010 42.590 4.280 ;
        RECT 43.430 0.010 43.510 4.280 ;
        RECT 44.350 0.010 44.430 4.280 ;
        RECT 45.270 0.010 45.350 4.280 ;
        RECT 46.190 0.010 46.270 4.280 ;
        RECT 47.110 0.010 47.190 4.280 ;
        RECT 48.030 0.010 48.110 4.280 ;
        RECT 48.950 0.010 49.030 4.280 ;
        RECT 49.870 0.010 49.950 4.280 ;
        RECT 50.790 0.010 50.870 4.280 ;
        RECT 51.710 0.010 51.790 4.280 ;
        RECT 52.630 0.010 52.710 4.280 ;
        RECT 53.550 0.010 53.630 4.280 ;
        RECT 54.470 0.010 54.550 4.280 ;
        RECT 55.390 0.010 55.470 4.280 ;
        RECT 56.310 0.010 56.390 4.280 ;
        RECT 57.230 0.010 57.310 4.280 ;
        RECT 58.150 0.010 58.230 4.280 ;
        RECT 59.070 0.010 59.150 4.280 ;
        RECT 59.990 0.010 60.070 4.280 ;
        RECT 60.910 0.010 60.990 4.280 ;
        RECT 61.830 0.010 61.910 4.280 ;
        RECT 62.750 0.010 62.830 4.280 ;
        RECT 63.670 0.010 63.750 4.280 ;
        RECT 64.590 0.010 64.670 4.280 ;
        RECT 65.510 0.010 65.590 4.280 ;
        RECT 66.430 0.010 66.510 4.280 ;
        RECT 67.350 0.010 67.430 4.280 ;
        RECT 68.270 0.010 68.350 4.280 ;
        RECT 69.190 0.010 69.270 4.280 ;
        RECT 70.110 0.010 70.190 4.280 ;
        RECT 71.030 0.010 71.110 4.280 ;
        RECT 71.950 0.010 72.030 4.280 ;
        RECT 72.870 0.010 72.950 4.280 ;
        RECT 73.790 0.010 73.870 4.280 ;
        RECT 74.710 0.010 74.790 4.280 ;
        RECT 75.630 0.010 75.710 4.280 ;
        RECT 76.550 0.010 76.630 4.280 ;
        RECT 77.470 0.010 77.550 4.280 ;
        RECT 78.390 0.010 78.470 4.280 ;
        RECT 79.310 0.010 79.390 4.280 ;
        RECT 80.230 0.010 80.310 4.280 ;
        RECT 81.150 0.010 81.230 4.280 ;
        RECT 82.070 0.010 82.150 4.280 ;
        RECT 82.990 0.010 83.070 4.280 ;
        RECT 83.910 0.010 83.990 4.280 ;
        RECT 84.830 0.010 84.910 4.280 ;
        RECT 85.750 0.010 85.830 4.280 ;
        RECT 86.670 0.010 86.750 4.280 ;
        RECT 87.590 0.010 87.670 4.280 ;
        RECT 88.510 0.010 88.590 4.280 ;
        RECT 89.430 0.010 89.510 4.280 ;
        RECT 90.350 0.010 90.430 4.280 ;
        RECT 91.270 0.010 91.350 4.280 ;
        RECT 92.190 0.010 92.270 4.280 ;
        RECT 93.110 0.010 93.190 4.280 ;
        RECT 94.030 0.010 94.110 4.280 ;
        RECT 94.950 0.010 95.030 4.280 ;
        RECT 95.870 0.010 95.950 4.280 ;
        RECT 96.790 0.010 96.870 4.280 ;
        RECT 97.710 0.010 97.790 4.280 ;
        RECT 98.630 0.010 98.710 4.280 ;
        RECT 99.550 0.010 99.630 4.280 ;
        RECT 100.470 0.010 199.910 4.280 ;
        RECT 200.750 0.010 201.750 4.280 ;
        RECT 202.590 0.010 203.590 4.280 ;
        RECT 204.430 0.010 205.430 4.280 ;
        RECT 206.270 0.010 207.270 4.280 ;
        RECT 208.110 0.010 209.110 4.280 ;
        RECT 209.950 0.010 210.950 4.280 ;
        RECT 211.790 0.010 212.790 4.280 ;
        RECT 213.630 0.010 400.010 4.280 ;
        RECT 400.850 0.010 401.850 4.280 ;
        RECT 402.690 0.010 403.690 4.280 ;
        RECT 404.530 0.010 405.530 4.280 ;
        RECT 406.370 0.010 474.210 4.280 ;
      LAYER met3 ;
        RECT 2.365 20.760 474.340 194.305 ;
        RECT 4.400 19.360 474.340 20.760 ;
        RECT 2.365 18.040 474.340 19.360 ;
        RECT 4.400 16.640 474.340 18.040 ;
        RECT 2.365 15.320 474.340 16.640 ;
        RECT 4.400 13.920 474.340 15.320 ;
        RECT 2.365 12.600 474.340 13.920 ;
        RECT 4.400 11.200 474.340 12.600 ;
        RECT 2.365 9.880 474.340 11.200 ;
        RECT 4.400 8.480 474.340 9.880 ;
        RECT 2.365 7.160 474.340 8.480 ;
        RECT 4.400 5.760 474.340 7.160 ;
        RECT 2.365 4.440 474.340 5.760 ;
        RECT 4.400 3.040 474.340 4.440 ;
        RECT 2.365 1.720 474.340 3.040 ;
        RECT 4.400 0.320 474.340 1.720 ;
        RECT 2.365 0.175 474.340 0.320 ;
      LAYER met4 ;
        RECT 12.255 188.320 325.385 194.305 ;
        RECT 12.255 11.735 18.940 188.320 ;
        RECT 24.740 11.735 68.940 188.320 ;
        RECT 74.740 11.735 118.940 188.320 ;
        RECT 124.740 11.735 168.940 188.320 ;
        RECT 174.740 11.735 218.940 188.320 ;
        RECT 224.740 11.735 268.940 188.320 ;
        RECT 274.740 11.735 318.940 188.320 ;
        RECT 324.740 11.735 325.385 188.320 ;
  END
END wb_host
MACRO sar_adc
  CLASS BLOCK ;
  FOREIGN sar_adc ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 300.000 ;
  PIN analog_dac_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 296.000 9.110 300.000 ;
    END
  END analog_dac_out
  PIN analog_din
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 296.000 8.190 300.000 ;
    END
  END analog_din
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.830 4.000 ;
    END
  END clk
  PIN pulse1m_mclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END pulse1m_mclk
  PIN reg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END reg_ack
  PIN reg_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END reg_addr[0]
  PIN reg_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END reg_addr[1]
  PIN reg_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END reg_addr[2]
  PIN reg_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END reg_addr[3]
  PIN reg_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END reg_addr[4]
  PIN reg_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END reg_addr[5]
  PIN reg_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END reg_addr[6]
  PIN reg_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END reg_addr[7]
  PIN reg_be[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END reg_be[0]
  PIN reg_be[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END reg_be[1]
  PIN reg_be[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 4.000 ;
    END
  END reg_be[2]
  PIN reg_be[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END reg_be[3]
  PIN reg_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END reg_cs
  PIN reg_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END reg_rdata[0]
  PIN reg_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END reg_rdata[10]
  PIN reg_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END reg_rdata[11]
  PIN reg_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END reg_rdata[12]
  PIN reg_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END reg_rdata[13]
  PIN reg_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END reg_rdata[14]
  PIN reg_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END reg_rdata[15]
  PIN reg_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END reg_rdata[16]
  PIN reg_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END reg_rdata[17]
  PIN reg_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END reg_rdata[18]
  PIN reg_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END reg_rdata[19]
  PIN reg_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END reg_rdata[1]
  PIN reg_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END reg_rdata[20]
  PIN reg_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END reg_rdata[21]
  PIN reg_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END reg_rdata[22]
  PIN reg_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END reg_rdata[23]
  PIN reg_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END reg_rdata[24]
  PIN reg_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END reg_rdata[25]
  PIN reg_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END reg_rdata[26]
  PIN reg_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END reg_rdata[27]
  PIN reg_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END reg_rdata[28]
  PIN reg_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END reg_rdata[29]
  PIN reg_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END reg_rdata[2]
  PIN reg_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END reg_rdata[30]
  PIN reg_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END reg_rdata[31]
  PIN reg_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END reg_rdata[3]
  PIN reg_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END reg_rdata[4]
  PIN reg_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END reg_rdata[5]
  PIN reg_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END reg_rdata[6]
  PIN reg_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END reg_rdata[7]
  PIN reg_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END reg_rdata[8]
  PIN reg_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END reg_rdata[9]
  PIN reg_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END reg_wdata[0]
  PIN reg_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END reg_wdata[10]
  PIN reg_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END reg_wdata[11]
  PIN reg_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END reg_wdata[12]
  PIN reg_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END reg_wdata[13]
  PIN reg_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END reg_wdata[14]
  PIN reg_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END reg_wdata[15]
  PIN reg_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END reg_wdata[16]
  PIN reg_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END reg_wdata[17]
  PIN reg_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END reg_wdata[18]
  PIN reg_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END reg_wdata[19]
  PIN reg_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END reg_wdata[1]
  PIN reg_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END reg_wdata[20]
  PIN reg_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END reg_wdata[21]
  PIN reg_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END reg_wdata[22]
  PIN reg_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END reg_wdata[23]
  PIN reg_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END reg_wdata[24]
  PIN reg_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END reg_wdata[25]
  PIN reg_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END reg_wdata[26]
  PIN reg_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END reg_wdata[27]
  PIN reg_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END reg_wdata[28]
  PIN reg_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END reg_wdata[29]
  PIN reg_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END reg_wdata[2]
  PIN reg_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END reg_wdata[30]
  PIN reg_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END reg_wdata[31]
  PIN reg_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END reg_wdata[3]
  PIN reg_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END reg_wdata[4]
  PIN reg_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END reg_wdata[5]
  PIN reg_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END reg_wdata[6]
  PIN reg_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END reg_wdata[7]
  PIN reg_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END reg_wdata[8]
  PIN reg_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END reg_wdata[9]
  PIN reg_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END reg_wr
  PIN reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END reset_n
  PIN sar2dac[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 296.000 7.270 300.000 ;
    END
  END sar2dac[0]
  PIN sar2dac[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 296.000 6.350 300.000 ;
    END
  END sar2dac[1]
  PIN sar2dac[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 296.000 5.430 300.000 ;
    END
  END sar2dac[2]
  PIN sar2dac[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 296.000 4.510 300.000 ;
    END
  END sar2dac[3]
  PIN sar2dac[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 296.000 3.590 300.000 ;
    END
  END sar2dac[4]
  PIN sar2dac[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 296.000 2.670 300.000 ;
    END
  END sar2dac[5]
  PIN sar2dac[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 296.000 1.750 300.000 ;
    END
  END sar2dac[6]
  PIN sar2dac[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 296.000 0.830 300.000 ;
    END
  END sar2dac[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 470.090 10.640 473.590 288.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 425.090 10.640 428.590 288.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 380.090 10.640 383.590 288.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 335.090 10.640 338.590 288.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 290.090 10.640 293.590 288.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 245.090 10.640 248.590 288.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 200.090 10.640 203.590 288.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 155.090 10.640 158.590 288.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 110.090 10.640 113.590 288.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 65.090 10.640 68.590 288.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.090 10.640 23.590 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 447.590 10.640 451.090 288.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 402.590 10.640 406.090 288.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 357.590 10.640 361.090 288.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 312.590 10.640 316.090 288.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 267.590 10.640 271.090 288.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 222.590 10.640 226.090 288.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 177.590 10.640 181.090 288.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 132.590 10.640 136.090 288.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 87.590 10.640 91.090 288.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 42.590 10.640 46.090 288.560 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 475.290 10.880 478.790 288.320 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 430.290 10.880 433.790 288.320 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 385.290 10.880 388.790 288.320 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 340.290 10.880 343.790 288.320 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 295.290 10.880 298.790 288.320 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 250.290 10.880 253.790 288.320 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 205.290 10.880 208.790 288.320 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 160.290 10.880 163.790 288.320 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 115.290 10.880 118.790 288.320 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 70.290 10.880 73.790 288.320 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 25.290 10.880 28.790 288.320 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 452.790 10.880 456.290 288.320 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 407.790 10.880 411.290 288.320 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 362.790 10.880 366.290 288.320 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 317.790 10.880 321.290 288.320 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 272.790 10.880 276.290 288.320 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 227.790 10.880 231.290 288.320 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 182.790 10.880 186.290 288.320 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 137.790 10.880 141.290 288.320 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 92.790 10.880 96.290 288.320 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 47.790 10.880 51.290 288.320 ;
    END
  END vssd2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 288.405 ;
      LAYER met1 ;
        RECT 0.530 6.840 494.040 288.560 ;
      LAYER met2 ;
        RECT 1.110 295.720 1.190 296.000 ;
        RECT 2.030 295.720 2.110 296.000 ;
        RECT 2.950 295.720 3.030 296.000 ;
        RECT 3.870 295.720 3.950 296.000 ;
        RECT 4.790 295.720 4.870 296.000 ;
        RECT 5.710 295.720 5.790 296.000 ;
        RECT 6.630 295.720 6.710 296.000 ;
        RECT 7.550 295.720 7.630 296.000 ;
        RECT 8.470 295.720 8.550 296.000 ;
        RECT 9.390 295.720 473.410 296.000 ;
        RECT 0.560 4.280 473.410 295.720 ;
        RECT 1.110 4.000 1.190 4.280 ;
        RECT 2.030 4.000 2.110 4.280 ;
        RECT 2.950 4.000 3.030 4.280 ;
        RECT 3.870 4.000 3.950 4.280 ;
        RECT 4.790 4.000 4.870 4.280 ;
        RECT 5.710 4.000 5.790 4.280 ;
        RECT 6.630 4.000 6.710 4.280 ;
        RECT 7.550 4.000 7.630 4.280 ;
        RECT 8.470 4.000 8.550 4.280 ;
        RECT 9.390 4.000 9.470 4.280 ;
        RECT 10.310 4.000 10.390 4.280 ;
        RECT 11.230 4.000 11.310 4.280 ;
        RECT 12.150 4.000 12.230 4.280 ;
        RECT 13.070 4.000 13.150 4.280 ;
        RECT 13.990 4.000 14.070 4.280 ;
        RECT 14.910 4.000 14.990 4.280 ;
        RECT 15.830 4.000 15.910 4.280 ;
        RECT 16.750 4.000 16.830 4.280 ;
        RECT 17.670 4.000 17.750 4.280 ;
        RECT 18.590 4.000 18.670 4.280 ;
        RECT 19.510 4.000 19.590 4.280 ;
        RECT 20.430 4.000 20.510 4.280 ;
        RECT 21.350 4.000 21.430 4.280 ;
        RECT 22.270 4.000 22.350 4.280 ;
        RECT 23.190 4.000 23.270 4.280 ;
        RECT 24.110 4.000 24.190 4.280 ;
        RECT 25.030 4.000 25.110 4.280 ;
        RECT 25.950 4.000 26.030 4.280 ;
        RECT 26.870 4.000 26.950 4.280 ;
        RECT 27.790 4.000 27.870 4.280 ;
        RECT 28.710 4.000 28.790 4.280 ;
        RECT 29.630 4.000 29.710 4.280 ;
        RECT 30.550 4.000 30.630 4.280 ;
        RECT 31.470 4.000 31.550 4.280 ;
        RECT 32.390 4.000 32.470 4.280 ;
        RECT 33.310 4.000 33.390 4.280 ;
        RECT 34.230 4.000 34.310 4.280 ;
        RECT 35.150 4.000 35.230 4.280 ;
        RECT 36.070 4.000 36.150 4.280 ;
        RECT 36.990 4.000 37.070 4.280 ;
        RECT 37.910 4.000 37.990 4.280 ;
        RECT 38.830 4.000 38.910 4.280 ;
        RECT 39.750 4.000 39.830 4.280 ;
        RECT 40.670 4.000 40.750 4.280 ;
        RECT 41.590 4.000 41.670 4.280 ;
        RECT 42.510 4.000 42.590 4.280 ;
        RECT 43.430 4.000 43.510 4.280 ;
        RECT 44.350 4.000 44.430 4.280 ;
        RECT 45.270 4.000 45.350 4.280 ;
        RECT 46.190 4.000 46.270 4.280 ;
        RECT 47.110 4.000 47.190 4.280 ;
        RECT 48.030 4.000 48.110 4.280 ;
        RECT 48.950 4.000 49.030 4.280 ;
        RECT 49.870 4.000 49.950 4.280 ;
        RECT 50.790 4.000 50.870 4.280 ;
        RECT 51.710 4.000 51.790 4.280 ;
        RECT 52.630 4.000 52.710 4.280 ;
        RECT 53.550 4.000 53.630 4.280 ;
        RECT 54.470 4.000 54.550 4.280 ;
        RECT 55.390 4.000 55.470 4.280 ;
        RECT 56.310 4.000 56.390 4.280 ;
        RECT 57.230 4.000 57.310 4.280 ;
        RECT 58.150 4.000 58.230 4.280 ;
        RECT 59.070 4.000 59.150 4.280 ;
        RECT 59.990 4.000 60.070 4.280 ;
        RECT 60.910 4.000 60.990 4.280 ;
        RECT 61.830 4.000 61.910 4.280 ;
        RECT 62.750 4.000 62.830 4.280 ;
        RECT 63.670 4.000 63.750 4.280 ;
        RECT 64.590 4.000 64.670 4.280 ;
        RECT 65.510 4.000 65.590 4.280 ;
        RECT 66.430 4.000 66.510 4.280 ;
        RECT 67.350 4.000 67.430 4.280 ;
        RECT 68.270 4.000 68.350 4.280 ;
        RECT 69.190 4.000 69.270 4.280 ;
        RECT 70.110 4.000 70.190 4.280 ;
        RECT 71.030 4.000 71.110 4.280 ;
        RECT 71.950 4.000 72.030 4.280 ;
        RECT 72.870 4.000 72.950 4.280 ;
        RECT 73.790 4.000 73.870 4.280 ;
        RECT 74.710 4.000 74.790 4.280 ;
        RECT 75.630 4.000 473.410 4.280 ;
      LAYER met3 ;
        RECT 1.445 10.715 473.590 288.485 ;
  END
END sar_adc
MACRO DAC_8BIT
  CLASS BLOCK ;
  FOREIGN DAC_8BIT ;
  ORIGIN 0.000 0.000 ;
  SIZE 499.220 BY 320.560 ;
  PIN d0
    PORT
      LAYER li1 ;
        RECT 106.460 19.395 106.760 25.600 ;
    END
    PORT
      LAYER met2 ;
        RECT 106.710 0.000 107.290 4.000 ;
    END
  END d0
  PIN d1
    PORT
      LAYER li1 ;
        RECT 121.850 19.960 122.150 26.270 ;
    END
    PORT
      LAYER met2 ;
        RECT 124.095 0.000 124.675 4.000 ;
    END
  END d1
  PIN d2
    PORT
      LAYER li1 ;
        RECT 138.550 20.880 138.850 27.510 ;
    END
    PORT
      LAYER met2 ;
        RECT 139.380 0.000 139.960 10.345 ;
    END
  END d2
  PIN d3
    PORT
      LAYER li1 ;
        RECT 155.520 21.790 155.820 28.980 ;
    END
    PORT
      LAYER met2 ;
        RECT 157.775 0.000 158.355 10.345 ;
    END
  END d3
  PIN d4
    PORT
      LAYER li1 ;
        RECT 171.730 23.100 172.030 30.410 ;
    END
    PORT
      LAYER met2 ;
        RECT 175.845 0.000 176.425 10.340 ;
    END
  END d4
  PIN d5
    PORT
      LAYER li1 ;
        RECT 189.040 23.410 189.340 48.150 ;
    END
    PORT
      LAYER met2 ;
        RECT 193.520 0.000 194.100 10.340 ;
    END
  END d5
  PIN d6
    PORT
      LAYER li1 ;
        RECT 215.460 24.380 215.790 31.770 ;
    END
    PORT
      LAYER met2 ;
        RECT 220.960 0.000 221.540 10.345 ;
    END
  END d6
  PIN x2_out_v
    PORT
      LAYER li1 ;
        RECT 480.860 155.910 481.070 158.160 ;
    END
  END x2_out_v
  PIN x1_out_v
    PORT
      LAYER li1 ;
        RECT 480.750 161.920 480.980 163.420 ;
    END
  END x1_out_v
  PIN out_v
    PORT
      LAYER li1 ;
        RECT 481.825 160.250 482.600 160.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 484.820 160.105 499.220 160.705 ;
    END
  END out_v
  PIN d7
    PORT
      LAYER li1 ;
        RECT 469.650 159.460 469.835 159.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 467.920 149.270 499.220 150.070 ;
    END
  END d7
  PIN inp1
    PORT
      LAYER li1 ;
        RECT 3.980 278.435 4.270 278.670 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.995 280.105 4.885 320.560 ;
    END
  END inp1
  PIN x2_vref1
    PORT
      LAYER li1 ;
        RECT 103.880 34.250 104.390 35.180 ;
    END
  END x2_vref1
  PIN x1_vref5
    PORT
      LAYER li1 ;
        RECT 103.000 36.230 103.510 37.100 ;
    END
  END x1_vref5
  PIN inp2
    PORT
      LAYER met2 ;
        RECT 339.785 0.000 340.365 10.275 ;
    END
  END inp2

  PIN gnd
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 55.030 281.005 60.350 320.560 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.185 279.130 19.505 320.560 ;
    END
  END vdd
  OBS
      LAYER li1 ;
        RECT 0.000 278.840 481.825 283.120 ;
        RECT 0.000 278.265 3.810 278.840 ;
        RECT 4.440 278.265 481.825 278.840 ;
        RECT 0.000 163.590 481.825 278.265 ;
        RECT 0.000 161.750 480.580 163.590 ;
        RECT 481.150 161.750 481.825 163.590 ;
        RECT 0.000 160.740 481.825 161.750 ;
        RECT 0.000 160.090 481.655 160.740 ;
        RECT 0.000 159.290 469.480 160.090 ;
        RECT 470.005 160.080 481.655 160.090 ;
        RECT 470.005 159.290 481.825 160.080 ;
        RECT 0.000 158.330 481.825 159.290 ;
        RECT 0.000 155.740 480.690 158.330 ;
        RECT 481.240 155.740 481.825 158.330 ;
        RECT 0.000 48.320 481.825 155.740 ;
        RECT 0.000 37.270 188.870 48.320 ;
        RECT 0.000 36.060 102.830 37.270 ;
        RECT 103.680 36.060 188.870 37.270 ;
        RECT 0.000 35.350 188.870 36.060 ;
        RECT 0.000 34.080 103.710 35.350 ;
        RECT 104.560 34.080 188.870 35.350 ;
        RECT 0.000 30.580 188.870 34.080 ;
        RECT 0.000 29.150 171.560 30.580 ;
        RECT 0.000 27.680 155.350 29.150 ;
        RECT 0.000 26.440 138.380 27.680 ;
        RECT 0.000 25.770 121.680 26.440 ;
        RECT 0.000 19.225 106.290 25.770 ;
        RECT 106.930 19.790 121.680 25.770 ;
        RECT 122.320 20.710 138.380 26.440 ;
        RECT 139.020 21.620 155.350 27.680 ;
        RECT 155.990 22.930 171.560 29.150 ;
        RECT 172.200 23.240 188.870 30.580 ;
        RECT 189.510 31.940 481.825 48.320 ;
        RECT 189.510 24.210 215.290 31.940 ;
        RECT 215.960 24.210 481.825 31.940 ;
        RECT 189.510 23.240 481.825 24.210 ;
        RECT 172.200 22.930 481.825 23.240 ;
        RECT 155.990 21.620 481.825 22.930 ;
        RECT 139.020 20.710 481.825 21.620 ;
        RECT 122.320 19.790 481.825 20.710 ;
        RECT 106.930 19.225 481.825 19.790 ;
        RECT 0.000 19.150 481.825 19.225 ;
      LAYER met1 ;
        RECT 3.125 10.265 483.290 282.230 ;
      LAYER met2 ;
        RECT 3.125 279.825 3.715 318.560 ;
        RECT 5.165 279.825 485.000 318.560 ;
        RECT 3.125 158.550 485.000 279.825 ;
        RECT 3.125 157.530 469.390 158.550 ;
        RECT 470.645 157.530 485.000 158.550 ;
        RECT 3.125 10.625 485.000 157.530 ;
        RECT 3.125 4.280 139.100 10.625 ;
        RECT 3.125 4.000 106.430 4.280 ;
        RECT 107.570 4.000 123.815 4.280 ;
        RECT 124.955 4.000 139.100 4.280 ;
        RECT 140.240 4.000 157.495 10.625 ;
        RECT 158.635 10.620 220.680 10.625 ;
        RECT 158.635 4.000 175.565 10.620 ;
        RECT 176.705 4.000 193.240 10.620 ;
        RECT 194.380 4.000 220.680 10.620 ;
        RECT 221.820 10.555 485.000 10.625 ;
        RECT 221.820 4.000 339.505 10.555 ;
        RECT 340.645 4.000 485.000 10.555 ;
      LAYER met3 ;
        RECT 10.220 161.105 497.080 282.315 ;
        RECT 10.220 159.705 484.420 161.105 ;
        RECT 10.220 150.470 497.080 159.705 ;
        RECT 10.220 148.870 467.520 150.470 ;
        RECT 10.220 44.630 497.080 148.870 ;
      LAYER met4 ;
        RECT 10.230 278.730 13.785 282.810 ;
        RECT 19.905 280.605 54.630 282.810 ;
        RECT 60.750 280.605 474.450 282.810 ;
        RECT 19.905 278.730 474.450 280.605 ;
        RECT 10.230 166.410 474.450 278.730 ;
        RECT 10.230 162.560 473.680 166.410 ;
        RECT 10.230 45.490 474.450 162.560 ;
  END
END DAC_8BIT
MACRO scr1_top_wb
  CLASS BLOCK ;
  FOREIGN scr1_top_wb ;
  ORIGIN 0.000 0.000 ;
  SIZE 1600.000 BY 1200.000 ;
  PIN core_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 0.720 1604.000 1.320 ;
    END
  END core_clk
  PIN cpu_rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 3.440 1604.000 4.040 ;
    END
  END cpu_rst_n
  PIN fuse_mhartid[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 70.080 1604.000 70.680 ;
    END
  END fuse_mhartid[0]
  PIN fuse_mhartid[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 56.480 1604.000 57.080 ;
    END
  END fuse_mhartid[10]
  PIN fuse_mhartid[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 55.120 1604.000 55.720 ;
    END
  END fuse_mhartid[11]
  PIN fuse_mhartid[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 53.760 1604.000 54.360 ;
    END
  END fuse_mhartid[12]
  PIN fuse_mhartid[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 52.400 1604.000 53.000 ;
    END
  END fuse_mhartid[13]
  PIN fuse_mhartid[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 51.040 1604.000 51.640 ;
    END
  END fuse_mhartid[14]
  PIN fuse_mhartid[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 49.680 1604.000 50.280 ;
    END
  END fuse_mhartid[15]
  PIN fuse_mhartid[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 48.320 1604.000 48.920 ;
    END
  END fuse_mhartid[16]
  PIN fuse_mhartid[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 46.960 1604.000 47.560 ;
    END
  END fuse_mhartid[17]
  PIN fuse_mhartid[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 45.600 1604.000 46.200 ;
    END
  END fuse_mhartid[18]
  PIN fuse_mhartid[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 44.240 1604.000 44.840 ;
    END
  END fuse_mhartid[19]
  PIN fuse_mhartid[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 68.720 1604.000 69.320 ;
    END
  END fuse_mhartid[1]
  PIN fuse_mhartid[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 42.880 1604.000 43.480 ;
    END
  END fuse_mhartid[20]
  PIN fuse_mhartid[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 41.520 1604.000 42.120 ;
    END
  END fuse_mhartid[21]
  PIN fuse_mhartid[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 40.160 1604.000 40.760 ;
    END
  END fuse_mhartid[22]
  PIN fuse_mhartid[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 38.800 1604.000 39.400 ;
    END
  END fuse_mhartid[23]
  PIN fuse_mhartid[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 37.440 1604.000 38.040 ;
    END
  END fuse_mhartid[24]
  PIN fuse_mhartid[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 36.080 1604.000 36.680 ;
    END
  END fuse_mhartid[25]
  PIN fuse_mhartid[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 34.720 1604.000 35.320 ;
    END
  END fuse_mhartid[26]
  PIN fuse_mhartid[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 33.360 1604.000 33.960 ;
    END
  END fuse_mhartid[27]
  PIN fuse_mhartid[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 32.000 1604.000 32.600 ;
    END
  END fuse_mhartid[28]
  PIN fuse_mhartid[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 30.640 1604.000 31.240 ;
    END
  END fuse_mhartid[29]
  PIN fuse_mhartid[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 67.360 1604.000 67.960 ;
    END
  END fuse_mhartid[2]
  PIN fuse_mhartid[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 29.280 1604.000 29.880 ;
    END
  END fuse_mhartid[30]
  PIN fuse_mhartid[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 27.920 1604.000 28.520 ;
    END
  END fuse_mhartid[31]
  PIN fuse_mhartid[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 66.000 1604.000 66.600 ;
    END
  END fuse_mhartid[3]
  PIN fuse_mhartid[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 64.640 1604.000 65.240 ;
    END
  END fuse_mhartid[4]
  PIN fuse_mhartid[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 63.280 1604.000 63.880 ;
    END
  END fuse_mhartid[5]
  PIN fuse_mhartid[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 61.920 1604.000 62.520 ;
    END
  END fuse_mhartid[6]
  PIN fuse_mhartid[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 60.560 1604.000 61.160 ;
    END
  END fuse_mhartid[7]
  PIN fuse_mhartid[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 59.200 1604.000 59.800 ;
    END
  END fuse_mhartid[8]
  PIN fuse_mhartid[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 57.840 1604.000 58.440 ;
    END
  END fuse_mhartid[9]
  PIN irq_lines[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 25.200 1604.000 25.800 ;
    END
  END irq_lines[0]
  PIN irq_lines[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 11.600 1604.000 12.200 ;
    END
  END irq_lines[10]
  PIN irq_lines[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 10.240 1604.000 10.840 ;
    END
  END irq_lines[11]
  PIN irq_lines[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 8.880 1604.000 9.480 ;
    END
  END irq_lines[12]
  PIN irq_lines[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 7.520 1604.000 8.120 ;
    END
  END irq_lines[13]
  PIN irq_lines[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 6.160 1604.000 6.760 ;
    END
  END irq_lines[14]
  PIN irq_lines[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 4.800 1604.000 5.400 ;
    END
  END irq_lines[15]
  PIN irq_lines[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 23.840 1604.000 24.440 ;
    END
  END irq_lines[1]
  PIN irq_lines[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 22.480 1604.000 23.080 ;
    END
  END irq_lines[2]
  PIN irq_lines[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 21.120 1604.000 21.720 ;
    END
  END irq_lines[3]
  PIN irq_lines[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 19.760 1604.000 20.360 ;
    END
  END irq_lines[4]
  PIN irq_lines[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 18.400 1604.000 19.000 ;
    END
  END irq_lines[5]
  PIN irq_lines[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 17.040 1604.000 17.640 ;
    END
  END irq_lines[6]
  PIN irq_lines[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 15.680 1604.000 16.280 ;
    END
  END irq_lines[7]
  PIN irq_lines[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 14.320 1604.000 14.920 ;
    END
  END irq_lines[8]
  PIN irq_lines[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 12.960 1604.000 13.560 ;
    END
  END irq_lines[9]
  PIN pwrup_rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 3.440 4.000 4.040 ;
    END
  END pwrup_rst_n
  PIN riscv_debug[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 -4.000 500.390 4.000 ;
    END
  END riscv_debug[0]
  PIN riscv_debug[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 -4.000 518.790 4.000 ;
    END
  END riscv_debug[10]
  PIN riscv_debug[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 -4.000 520.630 4.000 ;
    END
  END riscv_debug[11]
  PIN riscv_debug[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 -4.000 522.470 4.000 ;
    END
  END riscv_debug[12]
  PIN riscv_debug[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 -4.000 524.310 4.000 ;
    END
  END riscv_debug[13]
  PIN riscv_debug[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 -4.000 526.150 4.000 ;
    END
  END riscv_debug[14]
  PIN riscv_debug[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 -4.000 527.990 4.000 ;
    END
  END riscv_debug[15]
  PIN riscv_debug[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 -4.000 529.830 4.000 ;
    END
  END riscv_debug[16]
  PIN riscv_debug[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 -4.000 531.670 4.000 ;
    END
  END riscv_debug[17]
  PIN riscv_debug[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 -4.000 533.510 4.000 ;
    END
  END riscv_debug[18]
  PIN riscv_debug[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 -4.000 535.350 4.000 ;
    END
  END riscv_debug[19]
  PIN riscv_debug[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 -4.000 502.230 4.000 ;
    END
  END riscv_debug[1]
  PIN riscv_debug[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 -4.000 537.190 4.000 ;
    END
  END riscv_debug[20]
  PIN riscv_debug[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 -4.000 539.030 4.000 ;
    END
  END riscv_debug[21]
  PIN riscv_debug[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 -4.000 540.870 4.000 ;
    END
  END riscv_debug[22]
  PIN riscv_debug[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 -4.000 542.710 4.000 ;
    END
  END riscv_debug[23]
  PIN riscv_debug[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 -4.000 544.550 4.000 ;
    END
  END riscv_debug[24]
  PIN riscv_debug[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 -4.000 546.390 4.000 ;
    END
  END riscv_debug[25]
  PIN riscv_debug[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 -4.000 548.230 4.000 ;
    END
  END riscv_debug[26]
  PIN riscv_debug[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 -4.000 550.070 4.000 ;
    END
  END riscv_debug[27]
  PIN riscv_debug[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 -4.000 551.910 4.000 ;
    END
  END riscv_debug[28]
  PIN riscv_debug[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 -4.000 553.750 4.000 ;
    END
  END riscv_debug[29]
  PIN riscv_debug[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 -4.000 504.070 4.000 ;
    END
  END riscv_debug[2]
  PIN riscv_debug[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 -4.000 555.590 4.000 ;
    END
  END riscv_debug[30]
  PIN riscv_debug[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 -4.000 557.430 4.000 ;
    END
  END riscv_debug[31]
  PIN riscv_debug[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 -4.000 559.270 4.000 ;
    END
  END riscv_debug[32]
  PIN riscv_debug[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 -4.000 561.110 4.000 ;
    END
  END riscv_debug[33]
  PIN riscv_debug[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 -4.000 562.950 4.000 ;
    END
  END riscv_debug[34]
  PIN riscv_debug[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 -4.000 564.790 4.000 ;
    END
  END riscv_debug[35]
  PIN riscv_debug[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 -4.000 566.630 4.000 ;
    END
  END riscv_debug[36]
  PIN riscv_debug[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 -4.000 568.470 4.000 ;
    END
  END riscv_debug[37]
  PIN riscv_debug[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 -4.000 570.310 4.000 ;
    END
  END riscv_debug[38]
  PIN riscv_debug[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 -4.000 572.150 4.000 ;
    END
  END riscv_debug[39]
  PIN riscv_debug[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 -4.000 505.910 4.000 ;
    END
  END riscv_debug[3]
  PIN riscv_debug[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 -4.000 573.990 4.000 ;
    END
  END riscv_debug[40]
  PIN riscv_debug[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 -4.000 575.830 4.000 ;
    END
  END riscv_debug[41]
  PIN riscv_debug[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 -4.000 577.670 4.000 ;
    END
  END riscv_debug[42]
  PIN riscv_debug[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 -4.000 579.510 4.000 ;
    END
  END riscv_debug[43]
  PIN riscv_debug[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 -4.000 581.350 4.000 ;
    END
  END riscv_debug[44]
  PIN riscv_debug[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 -4.000 583.190 4.000 ;
    END
  END riscv_debug[45]
  PIN riscv_debug[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 -4.000 585.030 4.000 ;
    END
  END riscv_debug[46]
  PIN riscv_debug[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 -4.000 586.870 4.000 ;
    END
  END riscv_debug[47]
  PIN riscv_debug[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 -4.000 588.710 4.000 ;
    END
  END riscv_debug[48]
  PIN riscv_debug[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.270 -4.000 590.550 4.000 ;
    END
  END riscv_debug[49]
  PIN riscv_debug[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 -4.000 507.750 4.000 ;
    END
  END riscv_debug[4]
  PIN riscv_debug[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 -4.000 592.390 4.000 ;
    END
  END riscv_debug[50]
  PIN riscv_debug[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 -4.000 594.230 4.000 ;
    END
  END riscv_debug[51]
  PIN riscv_debug[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 -4.000 596.070 4.000 ;
    END
  END riscv_debug[52]
  PIN riscv_debug[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 -4.000 597.910 4.000 ;
    END
  END riscv_debug[53]
  PIN riscv_debug[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 -4.000 599.750 4.000 ;
    END
  END riscv_debug[54]
  PIN riscv_debug[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 -4.000 601.590 4.000 ;
    END
  END riscv_debug[55]
  PIN riscv_debug[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 -4.000 603.430 4.000 ;
    END
  END riscv_debug[56]
  PIN riscv_debug[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 -4.000 605.270 4.000 ;
    END
  END riscv_debug[57]
  PIN riscv_debug[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 -4.000 607.110 4.000 ;
    END
  END riscv_debug[58]
  PIN riscv_debug[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 -4.000 608.950 4.000 ;
    END
  END riscv_debug[59]
  PIN riscv_debug[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 -4.000 509.590 4.000 ;
    END
  END riscv_debug[5]
  PIN riscv_debug[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 -4.000 610.790 4.000 ;
    END
  END riscv_debug[60]
  PIN riscv_debug[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 -4.000 612.630 4.000 ;
    END
  END riscv_debug[61]
  PIN riscv_debug[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 -4.000 614.470 4.000 ;
    END
  END riscv_debug[62]
  PIN riscv_debug[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.030 -4.000 616.310 4.000 ;
    END
  END riscv_debug[63]
  PIN riscv_debug[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 -4.000 511.430 4.000 ;
    END
  END riscv_debug[6]
  PIN riscv_debug[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 -4.000 513.270 4.000 ;
    END
  END riscv_debug[7]
  PIN riscv_debug[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 -4.000 515.110 4.000 ;
    END
  END riscv_debug[8]
  PIN riscv_debug[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 -4.000 516.950 4.000 ;
    END
  END riscv_debug[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 4.800 4.000 5.400 ;
    END
  END rst_n
  PIN rtc_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 2.080 1604.000 2.680 ;
    END
  END rtc_clk
  PIN soft_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 26.560 1604.000 27.160 ;
    END
  END soft_irq
  PIN sram_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 425.720 1604.000 426.320 ;
    END
  END sram_addr0[0]
  PIN sram_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 423.000 1604.000 423.600 ;
    END
  END sram_addr0[1]
  PIN sram_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 420.280 1604.000 420.880 ;
    END
  END sram_addr0[2]
  PIN sram_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 417.560 1604.000 418.160 ;
    END
  END sram_addr0[3]
  PIN sram_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 414.840 1604.000 415.440 ;
    END
  END sram_addr0[4]
  PIN sram_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 412.120 1604.000 412.720 ;
    END
  END sram_addr0[5]
  PIN sram_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 409.400 1604.000 410.000 ;
    END
  END sram_addr0[6]
  PIN sram_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 406.680 1604.000 407.280 ;
    END
  END sram_addr0[7]
  PIN sram_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 403.960 1604.000 404.560 ;
    END
  END sram_addr0[8]
  PIN sram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 824.880 1604.000 825.480 ;
    END
  END sram_addr1[0]
  PIN sram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 822.160 1604.000 822.760 ;
    END
  END sram_addr1[1]
  PIN sram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 819.440 1604.000 820.040 ;
    END
  END sram_addr1[2]
  PIN sram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 816.720 1604.000 817.320 ;
    END
  END sram_addr1[3]
  PIN sram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 814.000 1604.000 814.600 ;
    END
  END sram_addr1[4]
  PIN sram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 811.280 1604.000 811.880 ;
    END
  END sram_addr1[5]
  PIN sram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 808.560 1604.000 809.160 ;
    END
  END sram_addr1[6]
  PIN sram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 805.840 1604.000 806.440 ;
    END
  END sram_addr1[7]
  PIN sram_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 803.120 1604.000 803.720 ;
    END
  END sram_addr1[8]
  PIN sram_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 401.240 1604.000 401.840 ;
    END
  END sram_csb0
  PIN sram_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 800.400 1604.000 801.000 ;
    END
  END sram_csb1
  PIN sram_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 384.920 1604.000 385.520 ;
    END
  END sram_din0[0]
  PIN sram_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 357.720 1604.000 358.320 ;
    END
  END sram_din0[10]
  PIN sram_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 355.000 1604.000 355.600 ;
    END
  END sram_din0[11]
  PIN sram_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 352.280 1604.000 352.880 ;
    END
  END sram_din0[12]
  PIN sram_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 349.560 1604.000 350.160 ;
    END
  END sram_din0[13]
  PIN sram_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 346.840 1604.000 347.440 ;
    END
  END sram_din0[14]
  PIN sram_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 344.120 1604.000 344.720 ;
    END
  END sram_din0[15]
  PIN sram_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 341.400 1604.000 342.000 ;
    END
  END sram_din0[16]
  PIN sram_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 338.680 1604.000 339.280 ;
    END
  END sram_din0[17]
  PIN sram_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 335.960 1604.000 336.560 ;
    END
  END sram_din0[18]
  PIN sram_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 333.240 1604.000 333.840 ;
    END
  END sram_din0[19]
  PIN sram_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 382.200 1604.000 382.800 ;
    END
  END sram_din0[1]
  PIN sram_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 330.520 1604.000 331.120 ;
    END
  END sram_din0[20]
  PIN sram_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 327.800 1604.000 328.400 ;
    END
  END sram_din0[21]
  PIN sram_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 325.080 1604.000 325.680 ;
    END
  END sram_din0[22]
  PIN sram_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 322.360 1604.000 322.960 ;
    END
  END sram_din0[23]
  PIN sram_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 319.640 1604.000 320.240 ;
    END
  END sram_din0[24]
  PIN sram_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 316.920 1604.000 317.520 ;
    END
  END sram_din0[25]
  PIN sram_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 314.200 1604.000 314.800 ;
    END
  END sram_din0[26]
  PIN sram_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 311.480 1604.000 312.080 ;
    END
  END sram_din0[27]
  PIN sram_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 308.760 1604.000 309.360 ;
    END
  END sram_din0[28]
  PIN sram_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 306.040 1604.000 306.640 ;
    END
  END sram_din0[29]
  PIN sram_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 379.480 1604.000 380.080 ;
    END
  END sram_din0[2]
  PIN sram_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 303.320 1604.000 303.920 ;
    END
  END sram_din0[30]
  PIN sram_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 300.600 1604.000 301.200 ;
    END
  END sram_din0[31]
  PIN sram_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 376.760 1604.000 377.360 ;
    END
  END sram_din0[3]
  PIN sram_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 374.040 1604.000 374.640 ;
    END
  END sram_din0[4]
  PIN sram_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 371.320 1604.000 371.920 ;
    END
  END sram_din0[5]
  PIN sram_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 368.600 1604.000 369.200 ;
    END
  END sram_din0[6]
  PIN sram_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 365.880 1604.000 366.480 ;
    END
  END sram_din0[7]
  PIN sram_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 363.160 1604.000 363.760 ;
    END
  END sram_din0[8]
  PIN sram_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 360.440 1604.000 361.040 ;
    END
  END sram_din0[9]
  PIN sram_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 284.960 1604.000 285.560 ;
    END
  END sram_dout0[0]
  PIN sram_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 257.760 1604.000 258.360 ;
    END
  END sram_dout0[10]
  PIN sram_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 255.040 1604.000 255.640 ;
    END
  END sram_dout0[11]
  PIN sram_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 252.320 1604.000 252.920 ;
    END
  END sram_dout0[12]
  PIN sram_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 249.600 1604.000 250.200 ;
    END
  END sram_dout0[13]
  PIN sram_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 246.880 1604.000 247.480 ;
    END
  END sram_dout0[14]
  PIN sram_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 244.160 1604.000 244.760 ;
    END
  END sram_dout0[15]
  PIN sram_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 241.440 1604.000 242.040 ;
    END
  END sram_dout0[16]
  PIN sram_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 238.720 1604.000 239.320 ;
    END
  END sram_dout0[17]
  PIN sram_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 236.000 1604.000 236.600 ;
    END
  END sram_dout0[18]
  PIN sram_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 233.280 1604.000 233.880 ;
    END
  END sram_dout0[19]
  PIN sram_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 282.240 1604.000 282.840 ;
    END
  END sram_dout0[1]
  PIN sram_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 230.560 1604.000 231.160 ;
    END
  END sram_dout0[20]
  PIN sram_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 227.840 1604.000 228.440 ;
    END
  END sram_dout0[21]
  PIN sram_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 225.120 1604.000 225.720 ;
    END
  END sram_dout0[22]
  PIN sram_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 222.400 1604.000 223.000 ;
    END
  END sram_dout0[23]
  PIN sram_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 219.680 1604.000 220.280 ;
    END
  END sram_dout0[24]
  PIN sram_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 216.960 1604.000 217.560 ;
    END
  END sram_dout0[25]
  PIN sram_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 214.240 1604.000 214.840 ;
    END
  END sram_dout0[26]
  PIN sram_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 211.520 1604.000 212.120 ;
    END
  END sram_dout0[27]
  PIN sram_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 208.800 1604.000 209.400 ;
    END
  END sram_dout0[28]
  PIN sram_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 206.080 1604.000 206.680 ;
    END
  END sram_dout0[29]
  PIN sram_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 279.520 1604.000 280.120 ;
    END
  END sram_dout0[2]
  PIN sram_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 203.360 1604.000 203.960 ;
    END
  END sram_dout0[30]
  PIN sram_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 200.640 1604.000 201.240 ;
    END
  END sram_dout0[31]
  PIN sram_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 276.800 1604.000 277.400 ;
    END
  END sram_dout0[3]
  PIN sram_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 274.080 1604.000 274.680 ;
    END
  END sram_dout0[4]
  PIN sram_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 271.360 1604.000 271.960 ;
    END
  END sram_dout0[5]
  PIN sram_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 268.640 1604.000 269.240 ;
    END
  END sram_dout0[6]
  PIN sram_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 265.920 1604.000 266.520 ;
    END
  END sram_dout0[7]
  PIN sram_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 263.200 1604.000 263.800 ;
    END
  END sram_dout0[8]
  PIN sram_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 260.480 1604.000 261.080 ;
    END
  END sram_dout0[9]
  PIN sram_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 911.920 1604.000 912.520 ;
    END
  END sram_dout1[0]
  PIN sram_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 884.720 1604.000 885.320 ;
    END
  END sram_dout1[10]
  PIN sram_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 882.000 1604.000 882.600 ;
    END
  END sram_dout1[11]
  PIN sram_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 879.280 1604.000 879.880 ;
    END
  END sram_dout1[12]
  PIN sram_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 876.560 1604.000 877.160 ;
    END
  END sram_dout1[13]
  PIN sram_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 873.840 1604.000 874.440 ;
    END
  END sram_dout1[14]
  PIN sram_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 871.120 1604.000 871.720 ;
    END
  END sram_dout1[15]
  PIN sram_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 868.400 1604.000 869.000 ;
    END
  END sram_dout1[16]
  PIN sram_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 865.680 1604.000 866.280 ;
    END
  END sram_dout1[17]
  PIN sram_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 862.960 1604.000 863.560 ;
    END
  END sram_dout1[18]
  PIN sram_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 860.240 1604.000 860.840 ;
    END
  END sram_dout1[19]
  PIN sram_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 909.200 1604.000 909.800 ;
    END
  END sram_dout1[1]
  PIN sram_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 857.520 1604.000 858.120 ;
    END
  END sram_dout1[20]
  PIN sram_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 854.800 1604.000 855.400 ;
    END
  END sram_dout1[21]
  PIN sram_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 852.080 1604.000 852.680 ;
    END
  END sram_dout1[22]
  PIN sram_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 849.360 1604.000 849.960 ;
    END
  END sram_dout1[23]
  PIN sram_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 846.640 1604.000 847.240 ;
    END
  END sram_dout1[24]
  PIN sram_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 843.920 1604.000 844.520 ;
    END
  END sram_dout1[25]
  PIN sram_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 841.200 1604.000 841.800 ;
    END
  END sram_dout1[26]
  PIN sram_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 838.480 1604.000 839.080 ;
    END
  END sram_dout1[27]
  PIN sram_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 835.760 1604.000 836.360 ;
    END
  END sram_dout1[28]
  PIN sram_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 833.040 1604.000 833.640 ;
    END
  END sram_dout1[29]
  PIN sram_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 906.480 1604.000 907.080 ;
    END
  END sram_dout1[2]
  PIN sram_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 830.320 1604.000 830.920 ;
    END
  END sram_dout1[30]
  PIN sram_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 827.600 1604.000 828.200 ;
    END
  END sram_dout1[31]
  PIN sram_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 903.760 1604.000 904.360 ;
    END
  END sram_dout1[3]
  PIN sram_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 901.040 1604.000 901.640 ;
    END
  END sram_dout1[4]
  PIN sram_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 898.320 1604.000 898.920 ;
    END
  END sram_dout1[5]
  PIN sram_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 895.600 1604.000 896.200 ;
    END
  END sram_dout1[6]
  PIN sram_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 892.880 1604.000 893.480 ;
    END
  END sram_dout1[7]
  PIN sram_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 890.160 1604.000 890.760 ;
    END
  END sram_dout1[8]
  PIN sram_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 887.440 1604.000 888.040 ;
    END
  END sram_dout1[9]
  PIN sram_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 398.520 1604.000 399.120 ;
    END
  END sram_web0
  PIN sram_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 395.800 1604.000 396.400 ;
    END
  END sram_wmask0[0]
  PIN sram_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 393.080 1604.000 393.680 ;
    END
  END sram_wmask0[1]
  PIN sram_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 390.360 1604.000 390.960 ;
    END
  END sram_wmask0[2]
  PIN sram_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 387.640 1604.000 388.240 ;
    END
  END sram_wmask0[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.340 10.640 23.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.340 10.640 123.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 220.340 10.640 223.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 320.340 10.640 323.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 420.340 10.640 423.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 520.340 10.640 523.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 620.340 10.640 623.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 720.340 10.640 723.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 820.340 10.640 823.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 920.340 10.640 923.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1020.340 10.640 1023.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1120.340 10.640 1123.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1220.340 10.640 1223.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1320.340 10.640 1323.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1420.340 10.640 1423.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1520.340 10.640 1523.340 1188.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 70.340 10.640 73.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 170.340 10.640 173.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 270.340 10.640 273.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 370.340 10.640 373.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 470.340 10.640 473.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 570.340 10.640 573.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 670.340 10.640 673.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 770.340 10.640 773.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 870.340 10.640 873.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 970.340 10.640 973.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1070.340 10.640 1073.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1170.340 10.640 1173.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1270.340 10.640 1273.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1370.340 10.640 1373.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1470.340 10.640 1473.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1570.340 10.640 1573.340 1188.880 ;
    END
  END vssd1
  PIN wb_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 0.720 4.000 1.320 ;
    END
  END wb_clk
  PIN wb_rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2.080 4.000 2.680 ;
    END
  END wb_rst_n
  PIN wbd_dmem_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 1196.000 594.230 1204.000 ;
    END
  END wbd_dmem_ack_i
  PIN wbd_dmem_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 1196.000 530.750 1204.000 ;
    END
  END wbd_dmem_adr_o[0]
  PIN wbd_dmem_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 1196.000 521.550 1204.000 ;
    END
  END wbd_dmem_adr_o[10]
  PIN wbd_dmem_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 1196.000 520.630 1204.000 ;
    END
  END wbd_dmem_adr_o[11]
  PIN wbd_dmem_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 1196.000 519.710 1204.000 ;
    END
  END wbd_dmem_adr_o[12]
  PIN wbd_dmem_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 1196.000 518.790 1204.000 ;
    END
  END wbd_dmem_adr_o[13]
  PIN wbd_dmem_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 1196.000 517.870 1204.000 ;
    END
  END wbd_dmem_adr_o[14]
  PIN wbd_dmem_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 1196.000 516.950 1204.000 ;
    END
  END wbd_dmem_adr_o[15]
  PIN wbd_dmem_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 1196.000 516.030 1204.000 ;
    END
  END wbd_dmem_adr_o[16]
  PIN wbd_dmem_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 1196.000 515.110 1204.000 ;
    END
  END wbd_dmem_adr_o[17]
  PIN wbd_dmem_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 1196.000 514.190 1204.000 ;
    END
  END wbd_dmem_adr_o[18]
  PIN wbd_dmem_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 1196.000 513.270 1204.000 ;
    END
  END wbd_dmem_adr_o[19]
  PIN wbd_dmem_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 1196.000 529.830 1204.000 ;
    END
  END wbd_dmem_adr_o[1]
  PIN wbd_dmem_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 1196.000 512.350 1204.000 ;
    END
  END wbd_dmem_adr_o[20]
  PIN wbd_dmem_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 1196.000 511.430 1204.000 ;
    END
  END wbd_dmem_adr_o[21]
  PIN wbd_dmem_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 1196.000 510.510 1204.000 ;
    END
  END wbd_dmem_adr_o[22]
  PIN wbd_dmem_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 1196.000 509.590 1204.000 ;
    END
  END wbd_dmem_adr_o[23]
  PIN wbd_dmem_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 1196.000 508.670 1204.000 ;
    END
  END wbd_dmem_adr_o[24]
  PIN wbd_dmem_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 1196.000 507.750 1204.000 ;
    END
  END wbd_dmem_adr_o[25]
  PIN wbd_dmem_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 1196.000 506.830 1204.000 ;
    END
  END wbd_dmem_adr_o[26]
  PIN wbd_dmem_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 1196.000 505.910 1204.000 ;
    END
  END wbd_dmem_adr_o[27]
  PIN wbd_dmem_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 1196.000 504.990 1204.000 ;
    END
  END wbd_dmem_adr_o[28]
  PIN wbd_dmem_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 1196.000 504.070 1204.000 ;
    END
  END wbd_dmem_adr_o[29]
  PIN wbd_dmem_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 1196.000 528.910 1204.000 ;
    END
  END wbd_dmem_adr_o[2]
  PIN wbd_dmem_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 1196.000 503.150 1204.000 ;
    END
  END wbd_dmem_adr_o[30]
  PIN wbd_dmem_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 1196.000 502.230 1204.000 ;
    END
  END wbd_dmem_adr_o[31]
  PIN wbd_dmem_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 1196.000 527.990 1204.000 ;
    END
  END wbd_dmem_adr_o[3]
  PIN wbd_dmem_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 1196.000 527.070 1204.000 ;
    END
  END wbd_dmem_adr_o[4]
  PIN wbd_dmem_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 1196.000 526.150 1204.000 ;
    END
  END wbd_dmem_adr_o[5]
  PIN wbd_dmem_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 1196.000 525.230 1204.000 ;
    END
  END wbd_dmem_adr_o[6]
  PIN wbd_dmem_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 1196.000 524.310 1204.000 ;
    END
  END wbd_dmem_adr_o[7]
  PIN wbd_dmem_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 1196.000 523.390 1204.000 ;
    END
  END wbd_dmem_adr_o[8]
  PIN wbd_dmem_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 1196.000 522.470 1204.000 ;
    END
  END wbd_dmem_adr_o[9]
  PIN wbd_dmem_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 1196.000 593.310 1204.000 ;
    END
  END wbd_dmem_dat_i[0]
  PIN wbd_dmem_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 1196.000 584.110 1204.000 ;
    END
  END wbd_dmem_dat_i[10]
  PIN wbd_dmem_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 1196.000 583.190 1204.000 ;
    END
  END wbd_dmem_dat_i[11]
  PIN wbd_dmem_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 1196.000 582.270 1204.000 ;
    END
  END wbd_dmem_dat_i[12]
  PIN wbd_dmem_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 1196.000 581.350 1204.000 ;
    END
  END wbd_dmem_dat_i[13]
  PIN wbd_dmem_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 1196.000 580.430 1204.000 ;
    END
  END wbd_dmem_dat_i[14]
  PIN wbd_dmem_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 1196.000 579.510 1204.000 ;
    END
  END wbd_dmem_dat_i[15]
  PIN wbd_dmem_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 1196.000 578.590 1204.000 ;
    END
  END wbd_dmem_dat_i[16]
  PIN wbd_dmem_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 1196.000 577.670 1204.000 ;
    END
  END wbd_dmem_dat_i[17]
  PIN wbd_dmem_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 1196.000 576.750 1204.000 ;
    END
  END wbd_dmem_dat_i[18]
  PIN wbd_dmem_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 1196.000 575.830 1204.000 ;
    END
  END wbd_dmem_dat_i[19]
  PIN wbd_dmem_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 1196.000 592.390 1204.000 ;
    END
  END wbd_dmem_dat_i[1]
  PIN wbd_dmem_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 1196.000 574.910 1204.000 ;
    END
  END wbd_dmem_dat_i[20]
  PIN wbd_dmem_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 1196.000 573.990 1204.000 ;
    END
  END wbd_dmem_dat_i[21]
  PIN wbd_dmem_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 1196.000 573.070 1204.000 ;
    END
  END wbd_dmem_dat_i[22]
  PIN wbd_dmem_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 1196.000 572.150 1204.000 ;
    END
  END wbd_dmem_dat_i[23]
  PIN wbd_dmem_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 1196.000 571.230 1204.000 ;
    END
  END wbd_dmem_dat_i[24]
  PIN wbd_dmem_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 1196.000 570.310 1204.000 ;
    END
  END wbd_dmem_dat_i[25]
  PIN wbd_dmem_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 1196.000 569.390 1204.000 ;
    END
  END wbd_dmem_dat_i[26]
  PIN wbd_dmem_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 1196.000 568.470 1204.000 ;
    END
  END wbd_dmem_dat_i[27]
  PIN wbd_dmem_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 1196.000 567.550 1204.000 ;
    END
  END wbd_dmem_dat_i[28]
  PIN wbd_dmem_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 1196.000 566.630 1204.000 ;
    END
  END wbd_dmem_dat_i[29]
  PIN wbd_dmem_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 1196.000 591.470 1204.000 ;
    END
  END wbd_dmem_dat_i[2]
  PIN wbd_dmem_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 1196.000 565.710 1204.000 ;
    END
  END wbd_dmem_dat_i[30]
  PIN wbd_dmem_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 1196.000 564.790 1204.000 ;
    END
  END wbd_dmem_dat_i[31]
  PIN wbd_dmem_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.270 1196.000 590.550 1204.000 ;
    END
  END wbd_dmem_dat_i[3]
  PIN wbd_dmem_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 1196.000 589.630 1204.000 ;
    END
  END wbd_dmem_dat_i[4]
  PIN wbd_dmem_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 1196.000 588.710 1204.000 ;
    END
  END wbd_dmem_dat_i[5]
  PIN wbd_dmem_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 1196.000 587.790 1204.000 ;
    END
  END wbd_dmem_dat_i[6]
  PIN wbd_dmem_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 1196.000 586.870 1204.000 ;
    END
  END wbd_dmem_dat_i[7]
  PIN wbd_dmem_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 1196.000 585.950 1204.000 ;
    END
  END wbd_dmem_dat_i[8]
  PIN wbd_dmem_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 1196.000 585.030 1204.000 ;
    END
  END wbd_dmem_dat_i[9]
  PIN wbd_dmem_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 1196.000 563.870 1204.000 ;
    END
  END wbd_dmem_dat_o[0]
  PIN wbd_dmem_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 1196.000 554.670 1204.000 ;
    END
  END wbd_dmem_dat_o[10]
  PIN wbd_dmem_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 1196.000 553.750 1204.000 ;
    END
  END wbd_dmem_dat_o[11]
  PIN wbd_dmem_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 1196.000 552.830 1204.000 ;
    END
  END wbd_dmem_dat_o[12]
  PIN wbd_dmem_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 1196.000 551.910 1204.000 ;
    END
  END wbd_dmem_dat_o[13]
  PIN wbd_dmem_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 1196.000 550.990 1204.000 ;
    END
  END wbd_dmem_dat_o[14]
  PIN wbd_dmem_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 1196.000 550.070 1204.000 ;
    END
  END wbd_dmem_dat_o[15]
  PIN wbd_dmem_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 1196.000 549.150 1204.000 ;
    END
  END wbd_dmem_dat_o[16]
  PIN wbd_dmem_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 1196.000 548.230 1204.000 ;
    END
  END wbd_dmem_dat_o[17]
  PIN wbd_dmem_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 1196.000 547.310 1204.000 ;
    END
  END wbd_dmem_dat_o[18]
  PIN wbd_dmem_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 1196.000 546.390 1204.000 ;
    END
  END wbd_dmem_dat_o[19]
  PIN wbd_dmem_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 1196.000 562.950 1204.000 ;
    END
  END wbd_dmem_dat_o[1]
  PIN wbd_dmem_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 1196.000 545.470 1204.000 ;
    END
  END wbd_dmem_dat_o[20]
  PIN wbd_dmem_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 1196.000 544.550 1204.000 ;
    END
  END wbd_dmem_dat_o[21]
  PIN wbd_dmem_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 1196.000 543.630 1204.000 ;
    END
  END wbd_dmem_dat_o[22]
  PIN wbd_dmem_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 1196.000 542.710 1204.000 ;
    END
  END wbd_dmem_dat_o[23]
  PIN wbd_dmem_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 1196.000 541.790 1204.000 ;
    END
  END wbd_dmem_dat_o[24]
  PIN wbd_dmem_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 1196.000 540.870 1204.000 ;
    END
  END wbd_dmem_dat_o[25]
  PIN wbd_dmem_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 1196.000 539.950 1204.000 ;
    END
  END wbd_dmem_dat_o[26]
  PIN wbd_dmem_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 1196.000 539.030 1204.000 ;
    END
  END wbd_dmem_dat_o[27]
  PIN wbd_dmem_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 1196.000 538.110 1204.000 ;
    END
  END wbd_dmem_dat_o[28]
  PIN wbd_dmem_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 1196.000 537.190 1204.000 ;
    END
  END wbd_dmem_dat_o[29]
  PIN wbd_dmem_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 1196.000 562.030 1204.000 ;
    END
  END wbd_dmem_dat_o[2]
  PIN wbd_dmem_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.990 1196.000 536.270 1204.000 ;
    END
  END wbd_dmem_dat_o[30]
  PIN wbd_dmem_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 1196.000 535.350 1204.000 ;
    END
  END wbd_dmem_dat_o[31]
  PIN wbd_dmem_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 1196.000 561.110 1204.000 ;
    END
  END wbd_dmem_dat_o[3]
  PIN wbd_dmem_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 1196.000 560.190 1204.000 ;
    END
  END wbd_dmem_dat_o[4]
  PIN wbd_dmem_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 1196.000 559.270 1204.000 ;
    END
  END wbd_dmem_dat_o[5]
  PIN wbd_dmem_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 1196.000 558.350 1204.000 ;
    END
  END wbd_dmem_dat_o[6]
  PIN wbd_dmem_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 1196.000 557.430 1204.000 ;
    END
  END wbd_dmem_dat_o[7]
  PIN wbd_dmem_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 1196.000 556.510 1204.000 ;
    END
  END wbd_dmem_dat_o[8]
  PIN wbd_dmem_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 1196.000 555.590 1204.000 ;
    END
  END wbd_dmem_dat_o[9]
  PIN wbd_dmem_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 1196.000 595.150 1204.000 ;
    END
  END wbd_dmem_err_i
  PIN wbd_dmem_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 1196.000 534.430 1204.000 ;
    END
  END wbd_dmem_sel_o[0]
  PIN wbd_dmem_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 1196.000 533.510 1204.000 ;
    END
  END wbd_dmem_sel_o[1]
  PIN wbd_dmem_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 1196.000 532.590 1204.000 ;
    END
  END wbd_dmem_sel_o[2]
  PIN wbd_dmem_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 1196.000 531.670 1204.000 ;
    END
  END wbd_dmem_sel_o[3]
  PIN wbd_dmem_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 1196.000 500.390 1204.000 ;
    END
  END wbd_dmem_stb_o
  PIN wbd_dmem_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 1196.000 501.310 1204.000 ;
    END
  END wbd_dmem_we_o
  PIN wbd_imem_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 1196.000 94.670 1204.000 ;
    END
  END wbd_imem_ack_i
  PIN wbd_imem_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 1196.000 31.190 1204.000 ;
    END
  END wbd_imem_adr_o[0]
  PIN wbd_imem_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 1196.000 21.990 1204.000 ;
    END
  END wbd_imem_adr_o[10]
  PIN wbd_imem_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 1196.000 21.070 1204.000 ;
    END
  END wbd_imem_adr_o[11]
  PIN wbd_imem_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 1196.000 20.150 1204.000 ;
    END
  END wbd_imem_adr_o[12]
  PIN wbd_imem_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 1196.000 19.230 1204.000 ;
    END
  END wbd_imem_adr_o[13]
  PIN wbd_imem_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 1196.000 18.310 1204.000 ;
    END
  END wbd_imem_adr_o[14]
  PIN wbd_imem_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 1196.000 17.390 1204.000 ;
    END
  END wbd_imem_adr_o[15]
  PIN wbd_imem_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 1196.000 16.470 1204.000 ;
    END
  END wbd_imem_adr_o[16]
  PIN wbd_imem_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 1196.000 15.550 1204.000 ;
    END
  END wbd_imem_adr_o[17]
  PIN wbd_imem_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 1196.000 14.630 1204.000 ;
    END
  END wbd_imem_adr_o[18]
  PIN wbd_imem_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 1196.000 13.710 1204.000 ;
    END
  END wbd_imem_adr_o[19]
  PIN wbd_imem_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 1196.000 30.270 1204.000 ;
    END
  END wbd_imem_adr_o[1]
  PIN wbd_imem_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 1196.000 12.790 1204.000 ;
    END
  END wbd_imem_adr_o[20]
  PIN wbd_imem_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 1196.000 11.870 1204.000 ;
    END
  END wbd_imem_adr_o[21]
  PIN wbd_imem_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 1196.000 10.950 1204.000 ;
    END
  END wbd_imem_adr_o[22]
  PIN wbd_imem_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 1196.000 10.030 1204.000 ;
    END
  END wbd_imem_adr_o[23]
  PIN wbd_imem_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 1196.000 9.110 1204.000 ;
    END
  END wbd_imem_adr_o[24]
  PIN wbd_imem_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 1196.000 8.190 1204.000 ;
    END
  END wbd_imem_adr_o[25]
  PIN wbd_imem_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 1196.000 7.270 1204.000 ;
    END
  END wbd_imem_adr_o[26]
  PIN wbd_imem_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 1196.000 6.350 1204.000 ;
    END
  END wbd_imem_adr_o[27]
  PIN wbd_imem_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 1196.000 5.430 1204.000 ;
    END
  END wbd_imem_adr_o[28]
  PIN wbd_imem_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 1196.000 4.510 1204.000 ;
    END
  END wbd_imem_adr_o[29]
  PIN wbd_imem_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 1196.000 29.350 1204.000 ;
    END
  END wbd_imem_adr_o[2]
  PIN wbd_imem_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 1196.000 3.590 1204.000 ;
    END
  END wbd_imem_adr_o[30]
  PIN wbd_imem_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 1196.000 2.670 1204.000 ;
    END
  END wbd_imem_adr_o[31]
  PIN wbd_imem_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 1196.000 28.430 1204.000 ;
    END
  END wbd_imem_adr_o[3]
  PIN wbd_imem_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 1196.000 27.510 1204.000 ;
    END
  END wbd_imem_adr_o[4]
  PIN wbd_imem_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 1196.000 26.590 1204.000 ;
    END
  END wbd_imem_adr_o[5]
  PIN wbd_imem_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 1196.000 25.670 1204.000 ;
    END
  END wbd_imem_adr_o[6]
  PIN wbd_imem_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 1196.000 24.750 1204.000 ;
    END
  END wbd_imem_adr_o[7]
  PIN wbd_imem_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 1196.000 23.830 1204.000 ;
    END
  END wbd_imem_adr_o[8]
  PIN wbd_imem_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 1196.000 22.910 1204.000 ;
    END
  END wbd_imem_adr_o[9]
  PIN wbd_imem_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 1196.000 93.750 1204.000 ;
    END
  END wbd_imem_dat_i[0]
  PIN wbd_imem_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 1196.000 84.550 1204.000 ;
    END
  END wbd_imem_dat_i[10]
  PIN wbd_imem_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 1196.000 83.630 1204.000 ;
    END
  END wbd_imem_dat_i[11]
  PIN wbd_imem_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 1196.000 82.710 1204.000 ;
    END
  END wbd_imem_dat_i[12]
  PIN wbd_imem_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 1196.000 81.790 1204.000 ;
    END
  END wbd_imem_dat_i[13]
  PIN wbd_imem_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 1196.000 80.870 1204.000 ;
    END
  END wbd_imem_dat_i[14]
  PIN wbd_imem_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 1196.000 79.950 1204.000 ;
    END
  END wbd_imem_dat_i[15]
  PIN wbd_imem_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 1196.000 79.030 1204.000 ;
    END
  END wbd_imem_dat_i[16]
  PIN wbd_imem_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 1196.000 78.110 1204.000 ;
    END
  END wbd_imem_dat_i[17]
  PIN wbd_imem_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 1196.000 77.190 1204.000 ;
    END
  END wbd_imem_dat_i[18]
  PIN wbd_imem_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 1196.000 76.270 1204.000 ;
    END
  END wbd_imem_dat_i[19]
  PIN wbd_imem_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 1196.000 92.830 1204.000 ;
    END
  END wbd_imem_dat_i[1]
  PIN wbd_imem_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 1196.000 75.350 1204.000 ;
    END
  END wbd_imem_dat_i[20]
  PIN wbd_imem_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 1196.000 74.430 1204.000 ;
    END
  END wbd_imem_dat_i[21]
  PIN wbd_imem_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 1196.000 73.510 1204.000 ;
    END
  END wbd_imem_dat_i[22]
  PIN wbd_imem_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 1196.000 72.590 1204.000 ;
    END
  END wbd_imem_dat_i[23]
  PIN wbd_imem_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 1196.000 71.670 1204.000 ;
    END
  END wbd_imem_dat_i[24]
  PIN wbd_imem_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 1196.000 70.750 1204.000 ;
    END
  END wbd_imem_dat_i[25]
  PIN wbd_imem_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 1196.000 69.830 1204.000 ;
    END
  END wbd_imem_dat_i[26]
  PIN wbd_imem_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 1196.000 68.910 1204.000 ;
    END
  END wbd_imem_dat_i[27]
  PIN wbd_imem_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 1196.000 67.990 1204.000 ;
    END
  END wbd_imem_dat_i[28]
  PIN wbd_imem_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 1196.000 67.070 1204.000 ;
    END
  END wbd_imem_dat_i[29]
  PIN wbd_imem_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 1196.000 91.910 1204.000 ;
    END
  END wbd_imem_dat_i[2]
  PIN wbd_imem_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 1196.000 66.150 1204.000 ;
    END
  END wbd_imem_dat_i[30]
  PIN wbd_imem_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 1196.000 65.230 1204.000 ;
    END
  END wbd_imem_dat_i[31]
  PIN wbd_imem_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 1196.000 90.990 1204.000 ;
    END
  END wbd_imem_dat_i[3]
  PIN wbd_imem_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 1196.000 90.070 1204.000 ;
    END
  END wbd_imem_dat_i[4]
  PIN wbd_imem_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 1196.000 89.150 1204.000 ;
    END
  END wbd_imem_dat_i[5]
  PIN wbd_imem_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 1196.000 88.230 1204.000 ;
    END
  END wbd_imem_dat_i[6]
  PIN wbd_imem_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 1196.000 87.310 1204.000 ;
    END
  END wbd_imem_dat_i[7]
  PIN wbd_imem_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 1196.000 86.390 1204.000 ;
    END
  END wbd_imem_dat_i[8]
  PIN wbd_imem_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 1196.000 85.470 1204.000 ;
    END
  END wbd_imem_dat_i[9]
  PIN wbd_imem_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 1196.000 64.310 1204.000 ;
    END
  END wbd_imem_dat_o[0]
  PIN wbd_imem_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 1196.000 55.110 1204.000 ;
    END
  END wbd_imem_dat_o[10]
  PIN wbd_imem_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 1196.000 54.190 1204.000 ;
    END
  END wbd_imem_dat_o[11]
  PIN wbd_imem_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 1196.000 53.270 1204.000 ;
    END
  END wbd_imem_dat_o[12]
  PIN wbd_imem_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 1196.000 52.350 1204.000 ;
    END
  END wbd_imem_dat_o[13]
  PIN wbd_imem_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 1196.000 51.430 1204.000 ;
    END
  END wbd_imem_dat_o[14]
  PIN wbd_imem_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 1196.000 50.510 1204.000 ;
    END
  END wbd_imem_dat_o[15]
  PIN wbd_imem_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 1196.000 49.590 1204.000 ;
    END
  END wbd_imem_dat_o[16]
  PIN wbd_imem_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 1196.000 48.670 1204.000 ;
    END
  END wbd_imem_dat_o[17]
  PIN wbd_imem_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 1196.000 47.750 1204.000 ;
    END
  END wbd_imem_dat_o[18]
  PIN wbd_imem_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 1196.000 46.830 1204.000 ;
    END
  END wbd_imem_dat_o[19]
  PIN wbd_imem_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 1196.000 63.390 1204.000 ;
    END
  END wbd_imem_dat_o[1]
  PIN wbd_imem_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 1196.000 45.910 1204.000 ;
    END
  END wbd_imem_dat_o[20]
  PIN wbd_imem_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 1196.000 44.990 1204.000 ;
    END
  END wbd_imem_dat_o[21]
  PIN wbd_imem_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 1196.000 44.070 1204.000 ;
    END
  END wbd_imem_dat_o[22]
  PIN wbd_imem_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 1196.000 43.150 1204.000 ;
    END
  END wbd_imem_dat_o[23]
  PIN wbd_imem_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 1196.000 42.230 1204.000 ;
    END
  END wbd_imem_dat_o[24]
  PIN wbd_imem_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 1196.000 41.310 1204.000 ;
    END
  END wbd_imem_dat_o[25]
  PIN wbd_imem_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 1196.000 40.390 1204.000 ;
    END
  END wbd_imem_dat_o[26]
  PIN wbd_imem_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 1196.000 39.470 1204.000 ;
    END
  END wbd_imem_dat_o[27]
  PIN wbd_imem_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 1196.000 38.550 1204.000 ;
    END
  END wbd_imem_dat_o[28]
  PIN wbd_imem_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 1196.000 37.630 1204.000 ;
    END
  END wbd_imem_dat_o[29]
  PIN wbd_imem_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 1196.000 62.470 1204.000 ;
    END
  END wbd_imem_dat_o[2]
  PIN wbd_imem_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 1196.000 36.710 1204.000 ;
    END
  END wbd_imem_dat_o[30]
  PIN wbd_imem_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 1196.000 35.790 1204.000 ;
    END
  END wbd_imem_dat_o[31]
  PIN wbd_imem_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 1196.000 61.550 1204.000 ;
    END
  END wbd_imem_dat_o[3]
  PIN wbd_imem_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 1196.000 60.630 1204.000 ;
    END
  END wbd_imem_dat_o[4]
  PIN wbd_imem_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 1196.000 59.710 1204.000 ;
    END
  END wbd_imem_dat_o[5]
  PIN wbd_imem_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 1196.000 58.790 1204.000 ;
    END
  END wbd_imem_dat_o[6]
  PIN wbd_imem_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 1196.000 57.870 1204.000 ;
    END
  END wbd_imem_dat_o[7]
  PIN wbd_imem_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 1196.000 56.950 1204.000 ;
    END
  END wbd_imem_dat_o[8]
  PIN wbd_imem_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 1196.000 56.030 1204.000 ;
    END
  END wbd_imem_dat_o[9]
  PIN wbd_imem_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 1196.000 95.590 1204.000 ;
    END
  END wbd_imem_err_i
  PIN wbd_imem_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 1196.000 34.870 1204.000 ;
    END
  END wbd_imem_sel_o[0]
  PIN wbd_imem_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 1196.000 33.950 1204.000 ;
    END
  END wbd_imem_sel_o[1]
  PIN wbd_imem_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 1196.000 33.030 1204.000 ;
    END
  END wbd_imem_sel_o[2]
  PIN wbd_imem_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 1196.000 32.110 1204.000 ;
    END
  END wbd_imem_sel_o[3]
  PIN wbd_imem_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 1196.000 0.830 1204.000 ;
    END
  END wbd_imem_stb_o
  PIN wbd_imem_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 1196.000 1.750 1204.000 ;
    END
  END wbd_imem_we_o
  OBS
      LAYER li1 ;
        RECT 5.520 2.465 1596.975 1195.695 ;
      LAYER met1 ;
        RECT 0.530 2.420 1597.035 1196.080 ;
      LAYER met2 ;
        RECT 1.110 1195.720 1.190 1196.110 ;
        RECT 2.030 1195.720 2.110 1196.110 ;
        RECT 2.950 1195.720 3.030 1196.110 ;
        RECT 3.870 1195.720 3.950 1196.110 ;
        RECT 4.790 1195.720 4.870 1196.110 ;
        RECT 5.710 1195.720 5.790 1196.110 ;
        RECT 6.630 1195.720 6.710 1196.110 ;
        RECT 7.550 1195.720 7.630 1196.110 ;
        RECT 8.470 1195.720 8.550 1196.110 ;
        RECT 9.390 1195.720 9.470 1196.110 ;
        RECT 10.310 1195.720 10.390 1196.110 ;
        RECT 11.230 1195.720 11.310 1196.110 ;
        RECT 12.150 1195.720 12.230 1196.110 ;
        RECT 13.070 1195.720 13.150 1196.110 ;
        RECT 13.990 1195.720 14.070 1196.110 ;
        RECT 14.910 1195.720 14.990 1196.110 ;
        RECT 15.830 1195.720 15.910 1196.110 ;
        RECT 16.750 1195.720 16.830 1196.110 ;
        RECT 17.670 1195.720 17.750 1196.110 ;
        RECT 18.590 1195.720 18.670 1196.110 ;
        RECT 19.510 1195.720 19.590 1196.110 ;
        RECT 20.430 1195.720 20.510 1196.110 ;
        RECT 21.350 1195.720 21.430 1196.110 ;
        RECT 22.270 1195.720 22.350 1196.110 ;
        RECT 23.190 1195.720 23.270 1196.110 ;
        RECT 24.110 1195.720 24.190 1196.110 ;
        RECT 25.030 1195.720 25.110 1196.110 ;
        RECT 25.950 1195.720 26.030 1196.110 ;
        RECT 26.870 1195.720 26.950 1196.110 ;
        RECT 27.790 1195.720 27.870 1196.110 ;
        RECT 28.710 1195.720 28.790 1196.110 ;
        RECT 29.630 1195.720 29.710 1196.110 ;
        RECT 30.550 1195.720 30.630 1196.110 ;
        RECT 31.470 1195.720 31.550 1196.110 ;
        RECT 32.390 1195.720 32.470 1196.110 ;
        RECT 33.310 1195.720 33.390 1196.110 ;
        RECT 34.230 1195.720 34.310 1196.110 ;
        RECT 35.150 1195.720 35.230 1196.110 ;
        RECT 36.070 1195.720 36.150 1196.110 ;
        RECT 36.990 1195.720 37.070 1196.110 ;
        RECT 37.910 1195.720 37.990 1196.110 ;
        RECT 38.830 1195.720 38.910 1196.110 ;
        RECT 39.750 1195.720 39.830 1196.110 ;
        RECT 40.670 1195.720 40.750 1196.110 ;
        RECT 41.590 1195.720 41.670 1196.110 ;
        RECT 42.510 1195.720 42.590 1196.110 ;
        RECT 43.430 1195.720 43.510 1196.110 ;
        RECT 44.350 1195.720 44.430 1196.110 ;
        RECT 45.270 1195.720 45.350 1196.110 ;
        RECT 46.190 1195.720 46.270 1196.110 ;
        RECT 47.110 1195.720 47.190 1196.110 ;
        RECT 48.030 1195.720 48.110 1196.110 ;
        RECT 48.950 1195.720 49.030 1196.110 ;
        RECT 49.870 1195.720 49.950 1196.110 ;
        RECT 50.790 1195.720 50.870 1196.110 ;
        RECT 51.710 1195.720 51.790 1196.110 ;
        RECT 52.630 1195.720 52.710 1196.110 ;
        RECT 53.550 1195.720 53.630 1196.110 ;
        RECT 54.470 1195.720 54.550 1196.110 ;
        RECT 55.390 1195.720 55.470 1196.110 ;
        RECT 56.310 1195.720 56.390 1196.110 ;
        RECT 57.230 1195.720 57.310 1196.110 ;
        RECT 58.150 1195.720 58.230 1196.110 ;
        RECT 59.070 1195.720 59.150 1196.110 ;
        RECT 59.990 1195.720 60.070 1196.110 ;
        RECT 60.910 1195.720 60.990 1196.110 ;
        RECT 61.830 1195.720 61.910 1196.110 ;
        RECT 62.750 1195.720 62.830 1196.110 ;
        RECT 63.670 1195.720 63.750 1196.110 ;
        RECT 64.590 1195.720 64.670 1196.110 ;
        RECT 65.510 1195.720 65.590 1196.110 ;
        RECT 66.430 1195.720 66.510 1196.110 ;
        RECT 67.350 1195.720 67.430 1196.110 ;
        RECT 68.270 1195.720 68.350 1196.110 ;
        RECT 69.190 1195.720 69.270 1196.110 ;
        RECT 70.110 1195.720 70.190 1196.110 ;
        RECT 71.030 1195.720 71.110 1196.110 ;
        RECT 71.950 1195.720 72.030 1196.110 ;
        RECT 72.870 1195.720 72.950 1196.110 ;
        RECT 73.790 1195.720 73.870 1196.110 ;
        RECT 74.710 1195.720 74.790 1196.110 ;
        RECT 75.630 1195.720 75.710 1196.110 ;
        RECT 76.550 1195.720 76.630 1196.110 ;
        RECT 77.470 1195.720 77.550 1196.110 ;
        RECT 78.390 1195.720 78.470 1196.110 ;
        RECT 79.310 1195.720 79.390 1196.110 ;
        RECT 80.230 1195.720 80.310 1196.110 ;
        RECT 81.150 1195.720 81.230 1196.110 ;
        RECT 82.070 1195.720 82.150 1196.110 ;
        RECT 82.990 1195.720 83.070 1196.110 ;
        RECT 83.910 1195.720 83.990 1196.110 ;
        RECT 84.830 1195.720 84.910 1196.110 ;
        RECT 85.750 1195.720 85.830 1196.110 ;
        RECT 86.670 1195.720 86.750 1196.110 ;
        RECT 87.590 1195.720 87.670 1196.110 ;
        RECT 88.510 1195.720 88.590 1196.110 ;
        RECT 89.430 1195.720 89.510 1196.110 ;
        RECT 90.350 1195.720 90.430 1196.110 ;
        RECT 91.270 1195.720 91.350 1196.110 ;
        RECT 92.190 1195.720 92.270 1196.110 ;
        RECT 93.110 1195.720 93.190 1196.110 ;
        RECT 94.030 1195.720 94.110 1196.110 ;
        RECT 94.950 1195.720 95.030 1196.110 ;
        RECT 95.870 1195.720 499.830 1196.110 ;
        RECT 500.670 1195.720 500.750 1196.110 ;
        RECT 501.590 1195.720 501.670 1196.110 ;
        RECT 502.510 1195.720 502.590 1196.110 ;
        RECT 503.430 1195.720 503.510 1196.110 ;
        RECT 504.350 1195.720 504.430 1196.110 ;
        RECT 505.270 1195.720 505.350 1196.110 ;
        RECT 506.190 1195.720 506.270 1196.110 ;
        RECT 507.110 1195.720 507.190 1196.110 ;
        RECT 508.030 1195.720 508.110 1196.110 ;
        RECT 508.950 1195.720 509.030 1196.110 ;
        RECT 509.870 1195.720 509.950 1196.110 ;
        RECT 510.790 1195.720 510.870 1196.110 ;
        RECT 511.710 1195.720 511.790 1196.110 ;
        RECT 512.630 1195.720 512.710 1196.110 ;
        RECT 513.550 1195.720 513.630 1196.110 ;
        RECT 514.470 1195.720 514.550 1196.110 ;
        RECT 515.390 1195.720 515.470 1196.110 ;
        RECT 516.310 1195.720 516.390 1196.110 ;
        RECT 517.230 1195.720 517.310 1196.110 ;
        RECT 518.150 1195.720 518.230 1196.110 ;
        RECT 519.070 1195.720 519.150 1196.110 ;
        RECT 519.990 1195.720 520.070 1196.110 ;
        RECT 520.910 1195.720 520.990 1196.110 ;
        RECT 521.830 1195.720 521.910 1196.110 ;
        RECT 522.750 1195.720 522.830 1196.110 ;
        RECT 523.670 1195.720 523.750 1196.110 ;
        RECT 524.590 1195.720 524.670 1196.110 ;
        RECT 525.510 1195.720 525.590 1196.110 ;
        RECT 526.430 1195.720 526.510 1196.110 ;
        RECT 527.350 1195.720 527.430 1196.110 ;
        RECT 528.270 1195.720 528.350 1196.110 ;
        RECT 529.190 1195.720 529.270 1196.110 ;
        RECT 530.110 1195.720 530.190 1196.110 ;
        RECT 531.030 1195.720 531.110 1196.110 ;
        RECT 531.950 1195.720 532.030 1196.110 ;
        RECT 532.870 1195.720 532.950 1196.110 ;
        RECT 533.790 1195.720 533.870 1196.110 ;
        RECT 534.710 1195.720 534.790 1196.110 ;
        RECT 535.630 1195.720 535.710 1196.110 ;
        RECT 536.550 1195.720 536.630 1196.110 ;
        RECT 537.470 1195.720 537.550 1196.110 ;
        RECT 538.390 1195.720 538.470 1196.110 ;
        RECT 539.310 1195.720 539.390 1196.110 ;
        RECT 540.230 1195.720 540.310 1196.110 ;
        RECT 541.150 1195.720 541.230 1196.110 ;
        RECT 542.070 1195.720 542.150 1196.110 ;
        RECT 542.990 1195.720 543.070 1196.110 ;
        RECT 543.910 1195.720 543.990 1196.110 ;
        RECT 544.830 1195.720 544.910 1196.110 ;
        RECT 545.750 1195.720 545.830 1196.110 ;
        RECT 546.670 1195.720 546.750 1196.110 ;
        RECT 547.590 1195.720 547.670 1196.110 ;
        RECT 548.510 1195.720 548.590 1196.110 ;
        RECT 549.430 1195.720 549.510 1196.110 ;
        RECT 550.350 1195.720 550.430 1196.110 ;
        RECT 551.270 1195.720 551.350 1196.110 ;
        RECT 552.190 1195.720 552.270 1196.110 ;
        RECT 553.110 1195.720 553.190 1196.110 ;
        RECT 554.030 1195.720 554.110 1196.110 ;
        RECT 554.950 1195.720 555.030 1196.110 ;
        RECT 555.870 1195.720 555.950 1196.110 ;
        RECT 556.790 1195.720 556.870 1196.110 ;
        RECT 557.710 1195.720 557.790 1196.110 ;
        RECT 558.630 1195.720 558.710 1196.110 ;
        RECT 559.550 1195.720 559.630 1196.110 ;
        RECT 560.470 1195.720 560.550 1196.110 ;
        RECT 561.390 1195.720 561.470 1196.110 ;
        RECT 562.310 1195.720 562.390 1196.110 ;
        RECT 563.230 1195.720 563.310 1196.110 ;
        RECT 564.150 1195.720 564.230 1196.110 ;
        RECT 565.070 1195.720 565.150 1196.110 ;
        RECT 565.990 1195.720 566.070 1196.110 ;
        RECT 566.910 1195.720 566.990 1196.110 ;
        RECT 567.830 1195.720 567.910 1196.110 ;
        RECT 568.750 1195.720 568.830 1196.110 ;
        RECT 569.670 1195.720 569.750 1196.110 ;
        RECT 570.590 1195.720 570.670 1196.110 ;
        RECT 571.510 1195.720 571.590 1196.110 ;
        RECT 572.430 1195.720 572.510 1196.110 ;
        RECT 573.350 1195.720 573.430 1196.110 ;
        RECT 574.270 1195.720 574.350 1196.110 ;
        RECT 575.190 1195.720 575.270 1196.110 ;
        RECT 576.110 1195.720 576.190 1196.110 ;
        RECT 577.030 1195.720 577.110 1196.110 ;
        RECT 577.950 1195.720 578.030 1196.110 ;
        RECT 578.870 1195.720 578.950 1196.110 ;
        RECT 579.790 1195.720 579.870 1196.110 ;
        RECT 580.710 1195.720 580.790 1196.110 ;
        RECT 581.630 1195.720 581.710 1196.110 ;
        RECT 582.550 1195.720 582.630 1196.110 ;
        RECT 583.470 1195.720 583.550 1196.110 ;
        RECT 584.390 1195.720 584.470 1196.110 ;
        RECT 585.310 1195.720 585.390 1196.110 ;
        RECT 586.230 1195.720 586.310 1196.110 ;
        RECT 587.150 1195.720 587.230 1196.110 ;
        RECT 588.070 1195.720 588.150 1196.110 ;
        RECT 588.990 1195.720 589.070 1196.110 ;
        RECT 589.910 1195.720 589.990 1196.110 ;
        RECT 590.830 1195.720 590.910 1196.110 ;
        RECT 591.750 1195.720 591.830 1196.110 ;
        RECT 592.670 1195.720 592.750 1196.110 ;
        RECT 593.590 1195.720 593.670 1196.110 ;
        RECT 594.510 1195.720 594.590 1196.110 ;
        RECT 595.430 1195.720 1595.650 1196.110 ;
        RECT 0.560 4.280 1595.650 1195.720 ;
        RECT 0.560 0.835 499.830 4.280 ;
        RECT 500.670 0.835 501.670 4.280 ;
        RECT 502.510 0.835 503.510 4.280 ;
        RECT 504.350 0.835 505.350 4.280 ;
        RECT 506.190 0.835 507.190 4.280 ;
        RECT 508.030 0.835 509.030 4.280 ;
        RECT 509.870 0.835 510.870 4.280 ;
        RECT 511.710 0.835 512.710 4.280 ;
        RECT 513.550 0.835 514.550 4.280 ;
        RECT 515.390 0.835 516.390 4.280 ;
        RECT 517.230 0.835 518.230 4.280 ;
        RECT 519.070 0.835 520.070 4.280 ;
        RECT 520.910 0.835 521.910 4.280 ;
        RECT 522.750 0.835 523.750 4.280 ;
        RECT 524.590 0.835 525.590 4.280 ;
        RECT 526.430 0.835 527.430 4.280 ;
        RECT 528.270 0.835 529.270 4.280 ;
        RECT 530.110 0.835 531.110 4.280 ;
        RECT 531.950 0.835 532.950 4.280 ;
        RECT 533.790 0.835 534.790 4.280 ;
        RECT 535.630 0.835 536.630 4.280 ;
        RECT 537.470 0.835 538.470 4.280 ;
        RECT 539.310 0.835 540.310 4.280 ;
        RECT 541.150 0.835 542.150 4.280 ;
        RECT 542.990 0.835 543.990 4.280 ;
        RECT 544.830 0.835 545.830 4.280 ;
        RECT 546.670 0.835 547.670 4.280 ;
        RECT 548.510 0.835 549.510 4.280 ;
        RECT 550.350 0.835 551.350 4.280 ;
        RECT 552.190 0.835 553.190 4.280 ;
        RECT 554.030 0.835 555.030 4.280 ;
        RECT 555.870 0.835 556.870 4.280 ;
        RECT 557.710 0.835 558.710 4.280 ;
        RECT 559.550 0.835 560.550 4.280 ;
        RECT 561.390 0.835 562.390 4.280 ;
        RECT 563.230 0.835 564.230 4.280 ;
        RECT 565.070 0.835 566.070 4.280 ;
        RECT 566.910 0.835 567.910 4.280 ;
        RECT 568.750 0.835 569.750 4.280 ;
        RECT 570.590 0.835 571.590 4.280 ;
        RECT 572.430 0.835 573.430 4.280 ;
        RECT 574.270 0.835 575.270 4.280 ;
        RECT 576.110 0.835 577.110 4.280 ;
        RECT 577.950 0.835 578.950 4.280 ;
        RECT 579.790 0.835 580.790 4.280 ;
        RECT 581.630 0.835 582.630 4.280 ;
        RECT 583.470 0.835 584.470 4.280 ;
        RECT 585.310 0.835 586.310 4.280 ;
        RECT 587.150 0.835 588.150 4.280 ;
        RECT 588.990 0.835 589.990 4.280 ;
        RECT 590.830 0.835 591.830 4.280 ;
        RECT 592.670 0.835 593.670 4.280 ;
        RECT 594.510 0.835 595.510 4.280 ;
        RECT 596.350 0.835 597.350 4.280 ;
        RECT 598.190 0.835 599.190 4.280 ;
        RECT 600.030 0.835 601.030 4.280 ;
        RECT 601.870 0.835 602.870 4.280 ;
        RECT 603.710 0.835 604.710 4.280 ;
        RECT 605.550 0.835 606.550 4.280 ;
        RECT 607.390 0.835 608.390 4.280 ;
        RECT 609.230 0.835 610.230 4.280 ;
        RECT 611.070 0.835 612.070 4.280 ;
        RECT 612.910 0.835 613.910 4.280 ;
        RECT 614.750 0.835 615.750 4.280 ;
        RECT 616.590 0.835 1595.650 4.280 ;
      LAYER met3 ;
        RECT 4.000 912.920 1596.000 1188.805 ;
        RECT 4.000 911.520 1595.600 912.920 ;
        RECT 4.000 910.200 1596.000 911.520 ;
        RECT 4.000 908.800 1595.600 910.200 ;
        RECT 4.000 907.480 1596.000 908.800 ;
        RECT 4.000 906.080 1595.600 907.480 ;
        RECT 4.000 904.760 1596.000 906.080 ;
        RECT 4.000 903.360 1595.600 904.760 ;
        RECT 4.000 902.040 1596.000 903.360 ;
        RECT 4.000 900.640 1595.600 902.040 ;
        RECT 4.000 899.320 1596.000 900.640 ;
        RECT 4.000 897.920 1595.600 899.320 ;
        RECT 4.000 896.600 1596.000 897.920 ;
        RECT 4.000 895.200 1595.600 896.600 ;
        RECT 4.000 893.880 1596.000 895.200 ;
        RECT 4.000 892.480 1595.600 893.880 ;
        RECT 4.000 891.160 1596.000 892.480 ;
        RECT 4.000 889.760 1595.600 891.160 ;
        RECT 4.000 888.440 1596.000 889.760 ;
        RECT 4.000 887.040 1595.600 888.440 ;
        RECT 4.000 885.720 1596.000 887.040 ;
        RECT 4.000 884.320 1595.600 885.720 ;
        RECT 4.000 883.000 1596.000 884.320 ;
        RECT 4.000 881.600 1595.600 883.000 ;
        RECT 4.000 880.280 1596.000 881.600 ;
        RECT 4.000 878.880 1595.600 880.280 ;
        RECT 4.000 877.560 1596.000 878.880 ;
        RECT 4.000 876.160 1595.600 877.560 ;
        RECT 4.000 874.840 1596.000 876.160 ;
        RECT 4.000 873.440 1595.600 874.840 ;
        RECT 4.000 872.120 1596.000 873.440 ;
        RECT 4.000 870.720 1595.600 872.120 ;
        RECT 4.000 869.400 1596.000 870.720 ;
        RECT 4.000 868.000 1595.600 869.400 ;
        RECT 4.000 866.680 1596.000 868.000 ;
        RECT 4.000 865.280 1595.600 866.680 ;
        RECT 4.000 863.960 1596.000 865.280 ;
        RECT 4.000 862.560 1595.600 863.960 ;
        RECT 4.000 861.240 1596.000 862.560 ;
        RECT 4.000 859.840 1595.600 861.240 ;
        RECT 4.000 858.520 1596.000 859.840 ;
        RECT 4.000 857.120 1595.600 858.520 ;
        RECT 4.000 855.800 1596.000 857.120 ;
        RECT 4.000 854.400 1595.600 855.800 ;
        RECT 4.000 853.080 1596.000 854.400 ;
        RECT 4.000 851.680 1595.600 853.080 ;
        RECT 4.000 850.360 1596.000 851.680 ;
        RECT 4.000 848.960 1595.600 850.360 ;
        RECT 4.000 847.640 1596.000 848.960 ;
        RECT 4.000 846.240 1595.600 847.640 ;
        RECT 4.000 844.920 1596.000 846.240 ;
        RECT 4.000 843.520 1595.600 844.920 ;
        RECT 4.000 842.200 1596.000 843.520 ;
        RECT 4.000 840.800 1595.600 842.200 ;
        RECT 4.000 839.480 1596.000 840.800 ;
        RECT 4.000 838.080 1595.600 839.480 ;
        RECT 4.000 836.760 1596.000 838.080 ;
        RECT 4.000 835.360 1595.600 836.760 ;
        RECT 4.000 834.040 1596.000 835.360 ;
        RECT 4.000 832.640 1595.600 834.040 ;
        RECT 4.000 831.320 1596.000 832.640 ;
        RECT 4.000 829.920 1595.600 831.320 ;
        RECT 4.000 828.600 1596.000 829.920 ;
        RECT 4.000 827.200 1595.600 828.600 ;
        RECT 4.000 825.880 1596.000 827.200 ;
        RECT 4.000 824.480 1595.600 825.880 ;
        RECT 4.000 823.160 1596.000 824.480 ;
        RECT 4.000 821.760 1595.600 823.160 ;
        RECT 4.000 820.440 1596.000 821.760 ;
        RECT 4.000 819.040 1595.600 820.440 ;
        RECT 4.000 817.720 1596.000 819.040 ;
        RECT 4.000 816.320 1595.600 817.720 ;
        RECT 4.000 815.000 1596.000 816.320 ;
        RECT 4.000 813.600 1595.600 815.000 ;
        RECT 4.000 812.280 1596.000 813.600 ;
        RECT 4.000 810.880 1595.600 812.280 ;
        RECT 4.000 809.560 1596.000 810.880 ;
        RECT 4.000 808.160 1595.600 809.560 ;
        RECT 4.000 806.840 1596.000 808.160 ;
        RECT 4.000 805.440 1595.600 806.840 ;
        RECT 4.000 804.120 1596.000 805.440 ;
        RECT 4.000 802.720 1595.600 804.120 ;
        RECT 4.000 801.400 1596.000 802.720 ;
        RECT 4.000 800.000 1595.600 801.400 ;
        RECT 4.000 426.720 1596.000 800.000 ;
        RECT 4.000 425.320 1595.600 426.720 ;
        RECT 4.000 424.000 1596.000 425.320 ;
        RECT 4.000 422.600 1595.600 424.000 ;
        RECT 4.000 421.280 1596.000 422.600 ;
        RECT 4.000 419.880 1595.600 421.280 ;
        RECT 4.000 418.560 1596.000 419.880 ;
        RECT 4.000 417.160 1595.600 418.560 ;
        RECT 4.000 415.840 1596.000 417.160 ;
        RECT 4.000 414.440 1595.600 415.840 ;
        RECT 4.000 413.120 1596.000 414.440 ;
        RECT 4.000 411.720 1595.600 413.120 ;
        RECT 4.000 410.400 1596.000 411.720 ;
        RECT 4.000 409.000 1595.600 410.400 ;
        RECT 4.000 407.680 1596.000 409.000 ;
        RECT 4.000 406.280 1595.600 407.680 ;
        RECT 4.000 404.960 1596.000 406.280 ;
        RECT 4.000 403.560 1595.600 404.960 ;
        RECT 4.000 402.240 1596.000 403.560 ;
        RECT 4.000 400.840 1595.600 402.240 ;
        RECT 4.000 399.520 1596.000 400.840 ;
        RECT 4.000 398.120 1595.600 399.520 ;
        RECT 4.000 396.800 1596.000 398.120 ;
        RECT 4.000 395.400 1595.600 396.800 ;
        RECT 4.000 394.080 1596.000 395.400 ;
        RECT 4.000 392.680 1595.600 394.080 ;
        RECT 4.000 391.360 1596.000 392.680 ;
        RECT 4.000 389.960 1595.600 391.360 ;
        RECT 4.000 388.640 1596.000 389.960 ;
        RECT 4.000 387.240 1595.600 388.640 ;
        RECT 4.000 385.920 1596.000 387.240 ;
        RECT 4.000 384.520 1595.600 385.920 ;
        RECT 4.000 383.200 1596.000 384.520 ;
        RECT 4.000 381.800 1595.600 383.200 ;
        RECT 4.000 380.480 1596.000 381.800 ;
        RECT 4.000 379.080 1595.600 380.480 ;
        RECT 4.000 377.760 1596.000 379.080 ;
        RECT 4.000 376.360 1595.600 377.760 ;
        RECT 4.000 375.040 1596.000 376.360 ;
        RECT 4.000 373.640 1595.600 375.040 ;
        RECT 4.000 372.320 1596.000 373.640 ;
        RECT 4.000 370.920 1595.600 372.320 ;
        RECT 4.000 369.600 1596.000 370.920 ;
        RECT 4.000 368.200 1595.600 369.600 ;
        RECT 4.000 366.880 1596.000 368.200 ;
        RECT 4.000 365.480 1595.600 366.880 ;
        RECT 4.000 364.160 1596.000 365.480 ;
        RECT 4.000 362.760 1595.600 364.160 ;
        RECT 4.000 361.440 1596.000 362.760 ;
        RECT 4.000 360.040 1595.600 361.440 ;
        RECT 4.000 358.720 1596.000 360.040 ;
        RECT 4.000 357.320 1595.600 358.720 ;
        RECT 4.000 356.000 1596.000 357.320 ;
        RECT 4.000 354.600 1595.600 356.000 ;
        RECT 4.000 353.280 1596.000 354.600 ;
        RECT 4.000 351.880 1595.600 353.280 ;
        RECT 4.000 350.560 1596.000 351.880 ;
        RECT 4.000 349.160 1595.600 350.560 ;
        RECT 4.000 347.840 1596.000 349.160 ;
        RECT 4.000 346.440 1595.600 347.840 ;
        RECT 4.000 345.120 1596.000 346.440 ;
        RECT 4.000 343.720 1595.600 345.120 ;
        RECT 4.000 342.400 1596.000 343.720 ;
        RECT 4.000 341.000 1595.600 342.400 ;
        RECT 4.000 339.680 1596.000 341.000 ;
        RECT 4.000 338.280 1595.600 339.680 ;
        RECT 4.000 336.960 1596.000 338.280 ;
        RECT 4.000 335.560 1595.600 336.960 ;
        RECT 4.000 334.240 1596.000 335.560 ;
        RECT 4.000 332.840 1595.600 334.240 ;
        RECT 4.000 331.520 1596.000 332.840 ;
        RECT 4.000 330.120 1595.600 331.520 ;
        RECT 4.000 328.800 1596.000 330.120 ;
        RECT 4.000 327.400 1595.600 328.800 ;
        RECT 4.000 326.080 1596.000 327.400 ;
        RECT 4.000 324.680 1595.600 326.080 ;
        RECT 4.000 323.360 1596.000 324.680 ;
        RECT 4.000 321.960 1595.600 323.360 ;
        RECT 4.000 320.640 1596.000 321.960 ;
        RECT 4.000 319.240 1595.600 320.640 ;
        RECT 4.000 317.920 1596.000 319.240 ;
        RECT 4.000 316.520 1595.600 317.920 ;
        RECT 4.000 315.200 1596.000 316.520 ;
        RECT 4.000 313.800 1595.600 315.200 ;
        RECT 4.000 312.480 1596.000 313.800 ;
        RECT 4.000 311.080 1595.600 312.480 ;
        RECT 4.000 309.760 1596.000 311.080 ;
        RECT 4.000 308.360 1595.600 309.760 ;
        RECT 4.000 307.040 1596.000 308.360 ;
        RECT 4.000 305.640 1595.600 307.040 ;
        RECT 4.000 304.320 1596.000 305.640 ;
        RECT 4.000 302.920 1595.600 304.320 ;
        RECT 4.000 301.600 1596.000 302.920 ;
        RECT 4.000 300.200 1595.600 301.600 ;
        RECT 4.000 285.960 1596.000 300.200 ;
        RECT 4.000 284.560 1595.600 285.960 ;
        RECT 4.000 283.240 1596.000 284.560 ;
        RECT 4.000 281.840 1595.600 283.240 ;
        RECT 4.000 280.520 1596.000 281.840 ;
        RECT 4.000 279.120 1595.600 280.520 ;
        RECT 4.000 277.800 1596.000 279.120 ;
        RECT 4.000 276.400 1595.600 277.800 ;
        RECT 4.000 275.080 1596.000 276.400 ;
        RECT 4.000 273.680 1595.600 275.080 ;
        RECT 4.000 272.360 1596.000 273.680 ;
        RECT 4.000 270.960 1595.600 272.360 ;
        RECT 4.000 269.640 1596.000 270.960 ;
        RECT 4.000 268.240 1595.600 269.640 ;
        RECT 4.000 266.920 1596.000 268.240 ;
        RECT 4.000 265.520 1595.600 266.920 ;
        RECT 4.000 264.200 1596.000 265.520 ;
        RECT 4.000 262.800 1595.600 264.200 ;
        RECT 4.000 261.480 1596.000 262.800 ;
        RECT 4.000 260.080 1595.600 261.480 ;
        RECT 4.000 258.760 1596.000 260.080 ;
        RECT 4.000 257.360 1595.600 258.760 ;
        RECT 4.000 256.040 1596.000 257.360 ;
        RECT 4.000 254.640 1595.600 256.040 ;
        RECT 4.000 253.320 1596.000 254.640 ;
        RECT 4.000 251.920 1595.600 253.320 ;
        RECT 4.000 250.600 1596.000 251.920 ;
        RECT 4.000 249.200 1595.600 250.600 ;
        RECT 4.000 247.880 1596.000 249.200 ;
        RECT 4.000 246.480 1595.600 247.880 ;
        RECT 4.000 245.160 1596.000 246.480 ;
        RECT 4.000 243.760 1595.600 245.160 ;
        RECT 4.000 242.440 1596.000 243.760 ;
        RECT 4.000 241.040 1595.600 242.440 ;
        RECT 4.000 239.720 1596.000 241.040 ;
        RECT 4.000 238.320 1595.600 239.720 ;
        RECT 4.000 237.000 1596.000 238.320 ;
        RECT 4.000 235.600 1595.600 237.000 ;
        RECT 4.000 234.280 1596.000 235.600 ;
        RECT 4.000 232.880 1595.600 234.280 ;
        RECT 4.000 231.560 1596.000 232.880 ;
        RECT 4.000 230.160 1595.600 231.560 ;
        RECT 4.000 228.840 1596.000 230.160 ;
        RECT 4.000 227.440 1595.600 228.840 ;
        RECT 4.000 226.120 1596.000 227.440 ;
        RECT 4.000 224.720 1595.600 226.120 ;
        RECT 4.000 223.400 1596.000 224.720 ;
        RECT 4.000 222.000 1595.600 223.400 ;
        RECT 4.000 220.680 1596.000 222.000 ;
        RECT 4.000 219.280 1595.600 220.680 ;
        RECT 4.000 217.960 1596.000 219.280 ;
        RECT 4.000 216.560 1595.600 217.960 ;
        RECT 4.000 215.240 1596.000 216.560 ;
        RECT 4.000 213.840 1595.600 215.240 ;
        RECT 4.000 212.520 1596.000 213.840 ;
        RECT 4.000 211.120 1595.600 212.520 ;
        RECT 4.000 209.800 1596.000 211.120 ;
        RECT 4.000 208.400 1595.600 209.800 ;
        RECT 4.000 207.080 1596.000 208.400 ;
        RECT 4.000 205.680 1595.600 207.080 ;
        RECT 4.000 204.360 1596.000 205.680 ;
        RECT 4.000 202.960 1595.600 204.360 ;
        RECT 4.000 201.640 1596.000 202.960 ;
        RECT 4.000 200.240 1595.600 201.640 ;
        RECT 4.000 71.080 1596.000 200.240 ;
        RECT 4.000 5.800 1595.600 71.080 ;
        RECT 4.400 0.855 1595.600 5.800 ;
      LAYER met4 ;
        RECT 376.575 12.415 419.940 1187.105 ;
        RECT 423.740 12.415 469.940 1187.105 ;
        RECT 473.740 12.415 519.940 1187.105 ;
        RECT 523.740 12.415 569.940 1187.105 ;
        RECT 573.740 12.415 619.940 1187.105 ;
        RECT 623.740 12.415 669.940 1187.105 ;
        RECT 673.740 12.415 719.940 1187.105 ;
        RECT 723.740 12.415 769.940 1187.105 ;
        RECT 773.740 12.415 819.940 1187.105 ;
        RECT 823.740 12.415 869.940 1187.105 ;
        RECT 873.740 12.415 919.940 1187.105 ;
        RECT 923.740 12.415 969.940 1187.105 ;
        RECT 973.740 12.415 1019.940 1187.105 ;
        RECT 1023.740 12.415 1069.940 1187.105 ;
        RECT 1073.740 12.415 1119.940 1187.105 ;
        RECT 1123.740 12.415 1169.940 1187.105 ;
        RECT 1173.740 12.415 1177.305 1187.105 ;
  END
END scr1_top_wb
MACRO sky130_sram_2kbyte_1rw1r_32x512_8
   CLASS BLOCK ;
   SIZE 683.1 BY 416.54 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  115.6 0.0 115.98 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  121.04 0.0 121.42 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  127.16 0.0 127.54 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  132.6 0.0 132.98 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  138.04 0.0 138.42 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  143.48 0.0 143.86 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  150.28 0.0 150.66 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  156.4 0.0 156.78 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  161.84 0.0 162.22 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  167.28 0.0 167.66 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  172.72 0.0 173.1 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  179.52 0.0 179.9 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  184.96 0.0 185.34 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  190.4 0.0 190.78 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  197.2 0.0 197.58 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  203.32 0.0 203.7 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  208.76 0.0 209.14 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  214.2 0.0 214.58 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  219.64 0.0 220.02 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  226.44 0.0 226.82 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  231.88 0.0 232.26 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  238.0 0.0 238.38 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  243.44 0.0 243.82 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  248.88 0.0 249.26 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  255.68 0.0 256.06 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  261.12 0.0 261.5 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  266.56 0.0 266.94 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  272.0 0.0 272.38 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  278.8 0.0 279.18 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  284.92 0.0 285.3 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  290.36 0.0 290.74 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  295.8 0.0 296.18 1.06 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  80.24 0.0 80.62 1.06 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  85.68 0.0 86.06 1.06 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 140.76 1.06 141.14 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 149.6 1.06 149.98 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 155.04 1.06 155.42 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 163.88 1.06 164.26 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 168.64 1.06 169.02 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 179.52 1.06 179.9 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 184.28 1.06 184.66 ;
      END
   END addr0[8]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  598.4 415.48 598.78 416.54 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  592.28 415.48 592.66 416.54 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 96.56 683.1 96.94 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 88.4 683.1 88.78 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 81.6 683.1 81.98 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 74.12 683.1 74.5 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 68.0 683.1 68.38 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  616.08 0.0 616.46 1.06 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  616.76 0.0 617.14 1.06 ;
      END
   END addr1[8]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 40.12 1.06 40.5 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 395.76 683.1 396.14 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 49.64 1.06 50.02 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 41.48 1.06 41.86 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  654.16 415.48 654.54 416.54 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  91.12 0.0 91.5 1.06 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  97.92 0.0 98.3 1.06 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  102.68 0.0 103.06 1.06 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  108.8 0.0 109.18 1.06 ;
      END
   END wmask0[3]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  141.44 0.0 141.82 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  153.68 0.0 154.06 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.96 0.0 168.34 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.2 0.0 180.58 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.44 0.0 192.82 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.36 0.0 205.74 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  217.6 0.0 217.98 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  229.84 0.0 230.22 1.06 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  241.4 0.0 241.78 1.06 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  255.0 0.0 255.38 1.06 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  267.92 0.0 268.3 1.06 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  280.16 0.0 280.54 1.06 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  292.4 0.0 292.78 1.06 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  304.64 0.0 305.02 1.06 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  317.56 0.0 317.94 1.06 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  329.8 0.0 330.18 1.06 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  341.36 0.0 341.74 1.06 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  354.96 0.0 355.34 1.06 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  367.2 0.0 367.58 1.06 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  379.44 0.0 379.82 1.06 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  392.36 0.0 392.74 1.06 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  404.6 0.0 404.98 1.06 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  417.52 0.0 417.9 1.06 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  429.76 0.0 430.14 1.06 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  442.68 0.0 443.06 1.06 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  454.92 0.0 455.3 1.06 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  467.16 0.0 467.54 1.06 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  479.4 0.0 479.78 1.06 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  492.32 0.0 492.7 1.06 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  504.56 0.0 504.94 1.06 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  516.8 0.0 517.18 1.06 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  529.72 0.0 530.1 1.06 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  143.48 415.48 143.86 416.54 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  155.04 415.48 155.42 416.54 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.28 415.48 167.66 416.54 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.88 415.48 181.26 416.54 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.44 415.48 192.82 416.54 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.36 415.48 205.74 416.54 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  217.6 415.48 217.98 416.54 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  230.52 415.48 230.9 416.54 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  242.76 415.48 243.14 416.54 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  255.68 415.48 256.06 416.54 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  267.92 415.48 268.3 416.54 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  280.84 415.48 281.22 416.54 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  292.4 415.48 292.78 416.54 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  304.64 415.48 305.02 416.54 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  318.24 415.48 318.62 416.54 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  330.48 415.48 330.86 416.54 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  342.72 415.48 343.1 416.54 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  354.96 415.48 355.34 416.54 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  367.88 415.48 368.26 416.54 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  379.44 415.48 379.82 416.54 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  393.04 415.48 393.42 416.54 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  405.28 415.48 405.66 416.54 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  417.52 415.48 417.9 416.54 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  429.76 415.48 430.14 416.54 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  442.0 415.48 442.38 416.54 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  454.92 415.48 455.3 416.54 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  467.84 415.48 468.22 416.54 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  480.08 415.48 480.46 416.54 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  492.32 415.48 492.7 416.54 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  505.24 415.48 505.62 416.54 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  516.8 415.48 517.18 416.54 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  530.4 415.48 530.78 416.54 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  4.76 4.76 6.5 411.78 ;
         LAYER met4 ;
         RECT  676.6 4.76 678.34 411.78 ;
         LAYER met3 ;
         RECT  4.76 410.04 678.34 411.78 ;
         LAYER met3 ;
         RECT  4.76 4.76 678.34 6.5 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  680.0 1.36 681.74 415.18 ;
         LAYER met4 ;
         RECT  1.36 1.36 3.1 415.18 ;
         LAYER met3 ;
         RECT  1.36 1.36 681.74 3.1 ;
         LAYER met3 ;
         RECT  1.36 413.44 681.74 415.18 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 682.48 415.92 ;
   LAYER  met2 ;
      RECT  0.62 0.62 682.48 415.92 ;
   LAYER  met3 ;
      RECT  1.66 140.16 682.48 141.74 ;
      RECT  0.62 141.74 1.66 149.0 ;
      RECT  0.62 150.58 1.66 154.44 ;
      RECT  0.62 156.02 1.66 163.28 ;
      RECT  0.62 164.86 1.66 168.04 ;
      RECT  0.62 169.62 1.66 178.92 ;
      RECT  0.62 180.5 1.66 183.68 ;
      RECT  1.66 95.96 681.44 97.54 ;
      RECT  1.66 97.54 681.44 140.16 ;
      RECT  681.44 97.54 682.48 140.16 ;
      RECT  681.44 89.38 682.48 95.96 ;
      RECT  681.44 82.58 682.48 87.8 ;
      RECT  681.44 75.1 682.48 81.0 ;
      RECT  681.44 68.98 682.48 73.52 ;
      RECT  1.66 141.74 681.44 395.16 ;
      RECT  1.66 395.16 681.44 396.74 ;
      RECT  681.44 141.74 682.48 395.16 ;
      RECT  0.62 50.62 1.66 140.16 ;
      RECT  0.62 42.46 1.66 49.04 ;
      RECT  1.66 396.74 4.16 409.44 ;
      RECT  1.66 409.44 4.16 412.38 ;
      RECT  4.16 396.74 678.94 409.44 ;
      RECT  678.94 396.74 681.44 409.44 ;
      RECT  678.94 409.44 681.44 412.38 ;
      RECT  1.66 4.16 4.16 7.1 ;
      RECT  1.66 7.1 4.16 95.96 ;
      RECT  4.16 7.1 678.94 95.96 ;
      RECT  678.94 4.16 681.44 7.1 ;
      RECT  678.94 7.1 681.44 95.96 ;
      RECT  681.44 0.62 682.34 0.76 ;
      RECT  681.44 3.7 682.34 67.4 ;
      RECT  682.34 0.62 682.48 0.76 ;
      RECT  682.34 0.76 682.48 3.7 ;
      RECT  682.34 3.7 682.48 67.4 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 39.52 ;
      RECT  0.76 0.62 1.66 0.76 ;
      RECT  0.76 3.7 1.66 39.52 ;
      RECT  1.66 0.62 4.16 0.76 ;
      RECT  1.66 3.7 4.16 4.16 ;
      RECT  4.16 0.62 678.94 0.76 ;
      RECT  4.16 3.7 678.94 4.16 ;
      RECT  678.94 0.62 681.44 0.76 ;
      RECT  678.94 3.7 681.44 4.16 ;
      RECT  0.62 185.26 0.76 412.84 ;
      RECT  0.62 412.84 0.76 415.78 ;
      RECT  0.62 415.78 0.76 415.92 ;
      RECT  0.76 185.26 1.66 412.84 ;
      RECT  0.76 415.78 1.66 415.92 ;
      RECT  681.44 396.74 682.34 412.84 ;
      RECT  681.44 415.78 682.34 415.92 ;
      RECT  682.34 396.74 682.48 412.84 ;
      RECT  682.34 412.84 682.48 415.78 ;
      RECT  682.34 415.78 682.48 415.92 ;
      RECT  1.66 412.38 4.16 412.84 ;
      RECT  1.66 415.78 4.16 415.92 ;
      RECT  4.16 412.38 678.94 412.84 ;
      RECT  4.16 415.78 678.94 415.92 ;
      RECT  678.94 412.38 681.44 412.84 ;
      RECT  678.94 415.78 681.44 415.92 ;
   LAYER  met4 ;
      RECT  115.0 1.66 116.58 415.92 ;
      RECT  116.58 0.62 120.44 1.66 ;
      RECT  122.02 0.62 126.56 1.66 ;
      RECT  128.14 0.62 132.0 1.66 ;
      RECT  133.58 0.62 137.44 1.66 ;
      RECT  144.46 0.62 149.68 1.66 ;
      RECT  157.38 0.62 161.24 1.66 ;
      RECT  162.82 0.62 166.68 1.66 ;
      RECT  173.7 0.62 178.92 1.66 ;
      RECT  185.94 0.62 189.8 1.66 ;
      RECT  198.18 0.62 202.72 1.66 ;
      RECT  209.74 0.62 213.6 1.66 ;
      RECT  220.62 0.62 225.84 1.66 ;
      RECT  232.86 0.62 237.4 1.66 ;
      RECT  244.42 0.62 248.28 1.66 ;
      RECT  256.66 0.62 260.52 1.66 ;
      RECT  262.1 0.62 265.96 1.66 ;
      RECT  272.98 0.62 278.2 1.66 ;
      RECT  285.9 0.62 289.76 1.66 ;
      RECT  81.22 0.62 85.08 1.66 ;
      RECT  116.58 1.66 597.8 414.88 ;
      RECT  597.8 1.66 599.38 414.88 ;
      RECT  593.26 414.88 597.8 415.92 ;
      RECT  599.38 414.88 653.56 415.92 ;
      RECT  86.66 0.62 90.52 1.66 ;
      RECT  92.1 0.62 97.32 1.66 ;
      RECT  98.9 0.62 102.08 1.66 ;
      RECT  103.66 0.62 108.2 1.66 ;
      RECT  109.78 0.62 115.0 1.66 ;
      RECT  139.02 0.62 140.84 1.66 ;
      RECT  142.42 0.62 142.88 1.66 ;
      RECT  151.26 0.62 153.08 1.66 ;
      RECT  154.66 0.62 155.8 1.66 ;
      RECT  168.94 0.62 172.12 1.66 ;
      RECT  181.18 0.62 184.36 1.66 ;
      RECT  191.38 0.62 191.84 1.66 ;
      RECT  193.42 0.62 196.6 1.66 ;
      RECT  204.3 0.62 204.76 1.66 ;
      RECT  206.34 0.62 208.16 1.66 ;
      RECT  215.18 0.62 217.0 1.66 ;
      RECT  218.58 0.62 219.04 1.66 ;
      RECT  227.42 0.62 229.24 1.66 ;
      RECT  230.82 0.62 231.28 1.66 ;
      RECT  238.98 0.62 240.8 1.66 ;
      RECT  242.38 0.62 242.84 1.66 ;
      RECT  249.86 0.62 254.4 1.66 ;
      RECT  268.9 0.62 271.4 1.66 ;
      RECT  281.14 0.62 284.32 1.66 ;
      RECT  291.34 0.62 291.8 1.66 ;
      RECT  293.38 0.62 295.2 1.66 ;
      RECT  296.78 0.62 304.04 1.66 ;
      RECT  305.62 0.62 316.96 1.66 ;
      RECT  318.54 0.62 329.2 1.66 ;
      RECT  330.78 0.62 340.76 1.66 ;
      RECT  342.34 0.62 354.36 1.66 ;
      RECT  355.94 0.62 366.6 1.66 ;
      RECT  368.18 0.62 378.84 1.66 ;
      RECT  380.42 0.62 391.76 1.66 ;
      RECT  393.34 0.62 404.0 1.66 ;
      RECT  405.58 0.62 416.92 1.66 ;
      RECT  418.5 0.62 429.16 1.66 ;
      RECT  430.74 0.62 442.08 1.66 ;
      RECT  443.66 0.62 454.32 1.66 ;
      RECT  455.9 0.62 466.56 1.66 ;
      RECT  468.14 0.62 478.8 1.66 ;
      RECT  480.38 0.62 491.72 1.66 ;
      RECT  493.3 0.62 503.96 1.66 ;
      RECT  505.54 0.62 516.2 1.66 ;
      RECT  517.78 0.62 529.12 1.66 ;
      RECT  530.7 0.62 615.48 1.66 ;
      RECT  116.58 414.88 142.88 415.92 ;
      RECT  144.46 414.88 154.44 415.92 ;
      RECT  156.02 414.88 166.68 415.92 ;
      RECT  168.26 414.88 180.28 415.92 ;
      RECT  181.86 414.88 191.84 415.92 ;
      RECT  193.42 414.88 204.76 415.92 ;
      RECT  206.34 414.88 217.0 415.92 ;
      RECT  218.58 414.88 229.92 415.92 ;
      RECT  231.5 414.88 242.16 415.92 ;
      RECT  243.74 414.88 255.08 415.92 ;
      RECT  256.66 414.88 267.32 415.92 ;
      RECT  268.9 414.88 280.24 415.92 ;
      RECT  281.82 414.88 291.8 415.92 ;
      RECT  293.38 414.88 304.04 415.92 ;
      RECT  305.62 414.88 317.64 415.92 ;
      RECT  319.22 414.88 329.88 415.92 ;
      RECT  331.46 414.88 342.12 415.92 ;
      RECT  343.7 414.88 354.36 415.92 ;
      RECT  355.94 414.88 367.28 415.92 ;
      RECT  368.86 414.88 378.84 415.92 ;
      RECT  380.42 414.88 392.44 415.92 ;
      RECT  394.02 414.88 404.68 415.92 ;
      RECT  406.26 414.88 416.92 415.92 ;
      RECT  418.5 414.88 429.16 415.92 ;
      RECT  430.74 414.88 441.4 415.92 ;
      RECT  442.98 414.88 454.32 415.92 ;
      RECT  455.9 414.88 467.24 415.92 ;
      RECT  468.82 414.88 479.48 415.92 ;
      RECT  481.06 414.88 491.72 415.92 ;
      RECT  493.3 414.88 504.64 415.92 ;
      RECT  506.22 414.88 516.2 415.92 ;
      RECT  517.78 414.88 529.8 415.92 ;
      RECT  531.38 414.88 591.68 415.92 ;
      RECT  4.16 1.66 7.1 4.16 ;
      RECT  4.16 412.38 7.1 415.92 ;
      RECT  7.1 1.66 115.0 4.16 ;
      RECT  7.1 4.16 115.0 412.38 ;
      RECT  7.1 412.38 115.0 415.92 ;
      RECT  599.38 1.66 676.0 4.16 ;
      RECT  599.38 4.16 676.0 412.38 ;
      RECT  599.38 412.38 676.0 414.88 ;
      RECT  676.0 1.66 678.94 4.16 ;
      RECT  676.0 412.38 678.94 414.88 ;
      RECT  617.74 0.62 679.4 0.76 ;
      RECT  617.74 0.76 679.4 1.66 ;
      RECT  679.4 0.62 682.34 0.76 ;
      RECT  682.34 0.62 682.48 0.76 ;
      RECT  682.34 0.76 682.48 1.66 ;
      RECT  655.14 414.88 679.4 415.78 ;
      RECT  655.14 415.78 679.4 415.92 ;
      RECT  679.4 415.78 682.34 415.92 ;
      RECT  682.34 414.88 682.48 415.78 ;
      RECT  682.34 415.78 682.48 415.92 ;
      RECT  678.94 1.66 679.4 4.16 ;
      RECT  682.34 1.66 682.48 4.16 ;
      RECT  678.94 4.16 679.4 412.38 ;
      RECT  682.34 4.16 682.48 412.38 ;
      RECT  678.94 412.38 679.4 414.88 ;
      RECT  682.34 412.38 682.48 414.88 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 1.66 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 79.64 0.76 ;
      RECT  3.7 0.76 79.64 1.66 ;
      RECT  0.62 1.66 0.76 4.16 ;
      RECT  3.7 1.66 4.16 4.16 ;
      RECT  0.62 4.16 0.76 412.38 ;
      RECT  3.7 4.16 4.16 412.38 ;
      RECT  0.62 412.38 0.76 415.78 ;
      RECT  0.62 415.78 0.76 415.92 ;
      RECT  0.76 415.78 3.7 415.92 ;
      RECT  3.7 412.38 4.16 415.78 ;
      RECT  3.7 415.78 4.16 415.92 ;
   END
END    sky130_sram_2kbyte_1rw1r_32x512_8
END LIBRARY